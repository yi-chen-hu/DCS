`define CYCLE_TIME 5.0

module PATTERN(
  // Input signals
	clk,
	rst_n,
    in_valid,
    in_cost,
  // Output signals
	out_valid,
    out_job,
	out_cost
);
//================================================================
// wire & registers 
//================================================================
output logic clk, rst_n, in_valid;
output logic [6:0] in_cost;
input out_valid;
input [3:0] out_job;
input [9:0] out_cost;

//================================================================
// clock
//================================================================
real	CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;

//================================================================
// parameters & integer
//================================================================
integer PATNUM = 250;
integer seed = 333;
integer i, j, k;
integer patcount;
integer gap;
integer input_file, output_file;

integer delay, out_cnt;
integer total_delay;
logic [9:0] golden_cost, design_cost[0:7];
logic [3:0] golden_job[0:7], design_job[0:7];
logic [6:0] golden_in [0:63];

integer SKIP = 0;
integer temp, s;
//================================================================
// initial
//================================================================
initial begin
	rst_n = 1'b1;
    in_valid = 1'b0;
	in_cost = 4'bx;
	total_delay = 0;

    input_file = $fopen("../00_TESTBED/input_TA.txt","r");
	output_file = $fopen("../00_TESTBED/output_TA.txt","r");
	skip_task;
	force clk = 0;
	reset_task;
	
	for(patcount=SKIP; patcount<PATNUM; patcount=patcount+1)
	begin	
		delay_task;	
		// $display("\033[33mPATTERN NO.%3d \033[m", patcount);
		input_task;
		ans_gen;
		wait_out_valid;
		check_ans;
		$display ("\033[0;32mPASS PATTERN NO.%3d, job: [ %1d, %1d, %1d, %1d, %1d, %1d, %1d, %1d], cost: %3d, Latency: %6d cycles\033[m", 
		patcount, 
		golden_job[0], golden_job[1], golden_job[2], golden_job[3], 
		golden_job[4], golden_job[5], golden_job[6], golden_job[7], golden_cost, delay);
	end

	YOU_PASS_task;
	$finish;
end

task reset_task ; begin
	#(2.5); rst_n = 0;

	#(50.0);
	if(out_valid !== 0 || out_job!==0 || out_cost!==0) begin
		fail;
		$display ("----------------------------------------------------------------------");
		$display ("                                FAIL!                                 ");
		$display ("              All output should be 0 after initial RESET              ");
		$display ("----------------------------------------------------------------------");
		#(100);
	    $finish ;
	end
	
	#(1.0); rst_n = 1 ;
	#(3.0); release clk;
end endtask


task delay_task; begin
	gap = $urandom_range(2,6);
	repeat(gap) @(negedge clk);
end endtask

task skip_task; begin
	for (s=0;s<SKIP;s=s+1) begin
		for (i=0;i<64;i=i+1)
			k = $fscanf(input_file, "%d", temp);
		for (i=0;i<9;i=i+1) 
			k = $fscanf(output_file, "%d", temp);
	end
end endtask

task input_task; begin
	in_valid = 1;
	for (i=0;i<64;i=i+1) begin
        k = $fscanf(input_file, "%d", in_cost);
		golden_in[i] = in_cost;
		@(negedge clk);
		check_out_while_input;
	end
	in_valid = 0;
	in_cost = 'dx;
	// $display("\033[34m     J1  J2  J3  J4  J5  J6  J7  J8\033[m",);
	// for (i=0;i<8;i=i+1) begin
		// $display("\033[34mW%1d: %3d %3d %3d %3d %3d %3d %3d %3d \033[m", 
		// i+1, golden_in[8*i], golden_in[8*i+1], golden_in[8*i+2], golden_in[8*i+3], golden_in[8*i+4], golden_in[8*i+5], golden_in[8*i+6], golden_in[8*i+7]);
	// end
end endtask

task ans_gen; begin
	for (i=0;i<8;i=i+1) 
		k = $fscanf(output_file, "%d", golden_job[i]);
	k = $fscanf(output_file, "%d", golden_cost);
end endtask

task check_out_while_input; begin
	if(in_valid===1 && out_valid!==0) begin
	fail;
	$display ("----------------------------------------------------------------------");
	$display ("                                FAIL!                                 ");
	$display ("                           Pattern No. %3d                            ",patcount);
	$display ("             out_valid should be 0 while in_valid is high             ");
	$display ("----------------------------------------------------------------------");
	#(100)
	$finish;
	end
end endtask

task wait_out_valid ; begin
	delay = 0;
	while(out_valid !== 1) begin
		@(negedge clk);
		delay = delay + 1;
		if(delay==400000) begin
			fail;
			$display ("----------------------------------------------------------------------");
			$display ("                                FAIL!                                 ");
			$display ("                           Pattern No. %3d                            ",patcount);
			$display ("            The execution latency are over 400,000 cycles             ");
			$display ("----------------------------------------------------------------------");
			#(100);
		    $finish ;
		end
	end
	total_delay = total_delay + delay;
end endtask

task check_ans; begin
	out_cnt = 0;
	for (i=0;i<8;i=i+1) begin	
		design_cost[i] = 'dx;
		design_job[i] = 'dx;
	end
	
	while (out_valid === 1) begin
		design_job[out_cnt] = out_job;
		design_cost[out_cnt] = out_cost;
		out_cnt = out_cnt + 1;
		if (out_cnt > 8) break;
		@(negedge clk);
	end
	
	if (out_cnt!=8) begin
		fail;
		$display ("----------------------------------------------------------------------");
		$display ("                                FAIL!                                 ");
		$display ("                           Pattern No. %3d                            ",patcount);
		$display ("              out_valid should be high only for 8 cycles              ");
		$display ("----------------------------------------------------------------------");
		#(100)
		$finish;
	end
	
	for (i=0;i<8;i=i+1) begin	
		if((design_job[i]!==golden_job[i]) || (design_cost[i]!=golden_cost)) begin
			fail;
			$display ("----------------------------------------------------------------------------------------------------");
			$display ("                                               FAIL!                                                ");
			$display ("                                          Pattern No. %3d                                           ",patcount);
			$display ("                                  J1  J2  J3  J4  J5  J6  J7  J8                                    ");
			for (j=0;j<8;j=j+1) begin
				if (golden_job[j]==1)
					$display ("                             W%1d: \033[94m%3d\033[m %3d %3d %3d %3d %3d %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==2)
					$display ("                             W%1d: %3d \033[94m%3d\033[m %3d %3d %3d %3d %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==3)
					$display ("                             W%1d: %3d %3d \033[94m%3d\033[m %3d %3d %3d %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==4)
					$display ("                             W%1d: %3d %3d %3d \033[94m%3d\033[m %3d %3d %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==5)
					$display ("                             W%1d: %3d %3d %3d %3d \033[94m%3d\033[m %3d %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==6)
					$display ("                             W%1d: %3d %3d %3d %3d %3d \033[94m%3d\033[m %3d %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==7)
					$display ("                             W%1d: %3d %3d %3d %3d %3d %3d \033[94m%3d\033[m %3d                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
				if (golden_job[j]==8)
					$display ("                             W%1d: %3d %3d %3d %3d %3d %3d %3d \033[94m%3d\033[m                                    ", 
					j+1, golden_in[8*j], golden_in[8*j+1], golden_in[8*j+2], golden_in[8*j+3], golden_in[8*j+4], golden_in[8*j+5], golden_in[8*j+6], golden_in[8*j+7]);
			end
			$display ("----------------------------------------------------------------------------------------------------");
			$display ("                   Your answer: job: [ %1d, %1d, %1d, %1d, %1d, %1d, %1d, %1d] cost: %3d                    ", 
			design_job[0], design_job[1], design_job[2], design_job[3], design_job[4], design_job[5], design_job[6], design_job[7], design_cost[i]);
			$display ("                   Gold answer: job: [ %1d, %1d, %1d, %1d, %1d, %1d, %1d, %1d] cost: %3d                    ", 
			golden_job[0], golden_job[1], golden_job[2], golden_job[3], golden_job[4], golden_job[5], golden_job[6], golden_job[7], golden_cost);
			$display ("-----------------------------------------------------------------------------------------------------");
			#(100)
			$finish;
		end
	end
	
	@(negedge clk);

end endtask

task YOU_PASS_task;begin
JohnCena;
// $display("\033[37m                                                                                                                                          ");        
// $display("\033[37m                                                                                \033[32m      :BBQvi.                                              ");        
// $display("\033[37m                                                              .i7ssrvs7         \033[32m     BBBBBBBBQi                                           ");        
// $display("\033[37m                        .:r7rrrr:::.        .::::::...   .i7vr:.      .B:       \033[32m    :BBBP :7BBBB.                                         ");        
// $display("\033[37m                      .Kv.........:rrvYr7v7rr:.....:rrirJr.   .rgBBBBg  Bi      \033[32m    BBBB     BBBB                                         ");        
// $display("\033[37m                     7Q  :rubEPUri:.       ..:irrii:..    :bBBBBBBBBBBB  B      \033[32m   iBBBv     BBBB       vBr                               ");        
// $display("\033[37m                    7B  BBBBBBBBBBBBBBB::BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB :R     \033[32m   BBBBBKrirBBBB.     :BBBBBB:                            ");        
// $display("\033[37m                   Jd .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: Bi    \033[32m  rBBBBBBBBBBBR.    .BBBM:BBB                             ");        
// $display("\033[37m                  uZ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B    \033[32m  BBBB   .::.      EBBBi :BBU                             ");        
// $display("\033[37m                 7B .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  B    \033[32m MBBBr           vBBBu   BBB.                             ");        
// $display("\033[37m                .B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: JJ   \033[32m i7PB          iBBBBB.  iBBB                              ");        
// $display("\033[37m                B. BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  Lu             \033[32m  vBBBBPBBBBPBBB7       .7QBB5i                ");        
// $display("\033[37m               Y1 KBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBi XBBBBBBBi :B            \033[32m :RBBB.  .rBBBBB.      rBBBBBBBB7              ");        
// $display("\033[37m              :B .BBBBBBBBBBBBBsRBBBBBBBBBBBrQBBBBB. UBBBRrBBBBBBr 1BBBBBBBBB  B.          \033[32m    .       BBBB       BBBB  :BBBB             ");        
// $display("\033[37m              Bi BBBBBBBBBBBBBi :BBBBBBBBBBE .BBK.  .  .   QBBBBBBBBBBBBBBBBBB  Bi         \033[32m           rBBBr       BBBB    BBBU            ");        
// $display("\033[37m             .B .BBBBBBBBBBBBBBQBBBBBBBBBBBB       \033[38;2;242;172;172mBBv \033[37m.LBBBBBBBBBBBBBBBBBBBBBB. B7.:ii:   \033[32m           vBBB        .BBBB   :7i.            ");        
// $display("\033[37m            .B  PBBBBBBBBBBBBBBBBBBBBBBBBBBBBbYQB. \033[38;2;242;172;172mBB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBB  Jr:::rK7 \033[32m             .7  BBB7   iBBBg                  ");        
// $display("\033[37m           7M  PBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBB..i   .   v1                  \033[32mdBBB.   5BBBr                 ");        
// $display("\033[37m          sZ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBB iD2BBQL.                 \033[32m ZBBBr  EBBBv     YBBBBQi     ");        
// $display("\033[37m  .7YYUSIX5 .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBBBY.:.      :B                 \033[32m  iBBBBBBBBD     BBBBBBBBB.   ");        
// $display("\033[37m LB.        ..BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB. \033[38;2;242;172;172mBB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBMBBB. BP17si                 \033[32m    :LBBBr      vBBBi  5BBB   ");        
// $display("\033[37m  KvJPBBB :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: \033[38;2;242;172;172mZB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBsiJr .i7ssr:                \033[32m          ...   :BBB:   BBBu  ");        
// $display("\033[37m i7ii:.   ::BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBj \033[38;2;242;172;172muBi \033[37mQBBBBBBBBBBBBBBBBBBBBBBBBi.ir      iB                \033[32m         .BBBi   BBBB   iMBu  ");        
// $display("\033[37mDB    .  vBdBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBg \033[38;2;242;172;172m7Bi \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBB rBrXPv.                \033[32m          BBBX   :BBBr        ");        
// $display("\033[37m :vQBBB. BQBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBQ \033[38;2;242;172;172miB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .L:ii::irrrrrrrr7jIr   \033[32m          .BBBv  :BBBQ        ");        
// $display("\033[37m :7:.   .. 5BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBr \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBB:            ..... ..YB. \033[32m           .BBBBBBBBB:        ");        
// $display("\033[37mBU  .:. BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mB7 \033[37mgBBBBBBBBBBBBBBBBBBBBBBBBBB. gBBBBBBBBBBBBBBBBBB. BL \033[32m             rBBBBB1.         ");        
// $display("\033[37m rY7iB: BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: \033[38;2;242;172;172mB7 \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBB. QBBBBBBBBBBBBBBBBBi  v5                                ");        
// $display("\033[37m     us EBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB \033[38;2;242;172;172mIr \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBgu7i.:BBBBBBBr Bu                                 ");        
// $display("\033[37m      B  7BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB.\033[38;2;242;172;172m:i \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBv:.  .. :::  .rr    rB                                  ");        
// $display("\033[37m      us  .BBBBBBBBBBBBBQLXBBBBBBBBBBBBBBBBBBBBBBBBq  .BBBBBBBBBBBBBBBBBBBBBBBBBv  :iJ7vri:::1Jr..isJYr                                   ");        
// $display("\033[37m      B  BBBBBBB  MBBBM      qBBBBBBBBBBBBBBBBBBBBBB: BBBBBBBBBBBBBBBBBBBBBBBBBB  B:           iir:                                       ");        
// $display("\033[37m     iB iBBBBBBBL       BBBP. :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  B.                                                       ");        
// $display("\033[37m     P: BBBBBBBBBBB5v7gBBBBBB  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: Br                                                        ");        
// $display("\033[37m     B  BBBs 7BBBBBBBBBBBBBB7 :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B                                                         ");        
// $display("\033[37m    .B :BBBB.  EBBBBBQBBBBBJ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB. B.                                                         ");        
// $display("\033[37m    ij qBBBBBg          ..  .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B                                                          ");        
// $display("\033[37m    UY QBBBBBBBBSUSPDQL...iBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBK EL                                                          ");        
// $display("\033[37m    B7 BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: B:                                                          ");        
// $display("\033[37m    B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBYrBB vBBBBBBBBBBBBBBBBBBBBBBBB. Ls                                                          ");        
// $display("\033[37m    B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBi_  /UBBBBBBBBBBBBBBBBBBBBBBBBB. :B:                                                        ");        
// $display("\033[37m   rM .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  ..IBBBBBBBBBBBBBBBBQBBBBBBBBBB  B                                                        ");        
// $display("\033[37m   B  BBBBBBBBBdZBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBPBBBBBBBBBBBBEji:..     sBBBBBBBr Br                                                       ");        
// $display("\033[37m  7B 7BBBBBBBr     .:vXQBBBBBBBBBBBBBBBBBBBBBBBBBQqui::..  ...i:i7777vi  BBBBBBr Bi                                                       ");        
// $display("\033[37m  Ki BBBBBBB  rY7vr:i....  .............:.....  ...:rii7vrr7r:..      7B  BBBBB  Bi                                                       ");        
// $display("\033[37m  B. BBBBBB  B:    .::ir77rrYLvvriiiiiiirvvY7rr77ri:..                 bU  iQBB:..rI                                                      ");        
// $display("\033[37m.S: 7BBBBP  B.                                                          vI7.  .:.  B.                                                     ");        
// $display("\033[37mB: ir:.   :B.                                                             :rvsUjUgU.                                                      ");        
// $display("\033[37mrMvrrirJKur                                                                                                                               \033[m");
$display ("----------------------------------------------------------------------------------------------------");
$display ("                                          Congratulations!                                          ");
$display ("                                    You have passed all patterns!                                   ");
$display ("                                    Total latency : %d cycles                                    ", total_delay);
$display ("----------------------------------------------------------------------------------------------------");

$finish;	
end endtask


task fail; begin
RickRoll;
// $display("\033[38;2;252;238;238m                                                                                                                                           ");      
// $display("\033[38;2;252;238;238m                                                                                                :L777777v7.                                ");
// $display("\033[31m  i:..::::::i.      :::::         ::::    .:::.       \033[38;2;252;238;238m                                       .vYr::::::::i7Lvi                             ");
// $display("\033[31m  BBBBBBBBBBBi     iBBBBBL       .BBBB    7BBB7       \033[38;2;252;238;238m                                      JL..\033[38;2;252;172;172m:r777v777i::\033[38;2;252;238;238m.ijL                           ");
// $display("\033[31m  BBBB.::::ir.     BBB:BBB.      .BBBv    iBBB:       \033[38;2;252;238;238m                                    :K: \033[38;2;252;172;172miv777rrrrr777v7:.\033[38;2;252;238;238m:J7                         ");
// $display("\033[31m  BBBQ            :BBY iBB7       BBB7    :BBB:       \033[38;2;252;238;238m                                   :d \033[38;2;252;172;172m.L7rrrrrrrrrrrrr77v: \033[38;2;252;238;238miI.                       ");
// $display("\033[31m  BBBB            BBB. .BBB.      BBB7    :BBB:       \033[38;2;252;238;238m                                  .B \033[38;2;252;172;172m.L7rrrrrrrrrrrrrrrrr7v..\033[38;2;252;238;238mBr                      ");
// $display("\033[31m  BBBB:r7vvj:    :BBB   gBBs      BBB7    :BBB:       \033[38;2;252;238;238m                                  S:\033[38;2;252;172;172m v7rrrrrrrrrrrrrrrrrrr7v. \033[38;2;252;238;238mB:                     ");
// $display("\033[31m  BBBBBBBBBB7    BBB:   .BBB.     BBB7    :BBB:       \033[38;2;252;238;238m                                 .D \033[38;2;252;172;172mi7rrrrrrr777rrrrrrrrrrr7v. \033[38;2;252;238;238mB.                    ");
// $display("\033[31m  BBBB    ..    iBBBBBBBBBBBP     BBB7    :BBB:       \033[38;2;252;238;238m                                 rv\033[38;2;252;172;172m v7rrrrrr7rirv7rrrrrrrrrr7v \033[38;2;252;238;238m:I                    ");
// $display("\033[31m  BBBB          BBBBi7vviQBBB.    BBB7    :BBB.       \033[38;2;252;238;238m                                 2i\033[38;2;252;172;172m.v7rrrrrr7i  :v7rrrrrrrrrrvi \033[38;2;252;238;238mB:                   ");
// $display("\033[31m  BBBB         rBBB.      BBBQ   .BBBv    iBBB2ir777L7\033[38;2;252;238;238m                                 2i.\033[38;2;252;172;172mv7rrrrrr7v \033[38;2;252;238;238m:..\033[38;2;252;172;172mv7rrrrrrrrr77 \033[38;2;252;238;238mrX                   ");
// $display("\033[31m .BBBB        :BBBB       BBBB7  .BBBB    7BBBBBBBBBBB\033[38;2;252;238;238m                                 Yv \033[38;2;252;172;172mv7rrrrrrrv.\033[38;2;252;238;238m.B \033[38;2;252;172;172m.vrrrrrrrrrrL.\033[38;2;252;238;238m:5                   ");
// $display("\033[31m  . ..        ....         ...:   ....    ..   .......\033[38;2;252;238;238m                                 .q \033[38;2;252;172;172mr7rrrrrrr7i \033[38;2;252;238;238mPv \033[38;2;252;172;172mi7rrrrrrrrrv.\033[38;2;252;238;238m:S                   ");
// $display("\033[38;2;252;238;238m                                                                                        Lr \033[38;2;252;172;172m77rrrrrr77 \033[38;2;252;238;238m:B. \033[38;2;252;172;172mv7rrrrrrrrv.\033[38;2;252;238;238m:S                   ");
// $display("\033[38;2;252;238;238m                                                                                         B: \033[38;2;252;172;172m7v7rrrrrv. \033[38;2;252;238;238mBY \033[38;2;252;172;172mi7rrrrrrr7v \033[38;2;252;238;238miK                   ");
// $display("\033[38;2;252;238;238m                                                                              .::rriii7rir7. \033[38;2;252;172;172m.r77777vi \033[38;2;252;238;238m7B  \033[38;2;252;172;172mvrrrrrrr7r \033[38;2;252;238;238m2r                   ");
// $display("\033[38;2;252;238;238m                                                                       .:rr7rri::......    .     \033[38;2;252;172;172m.:i7s \033[38;2;252;238;238m.B. \033[38;2;252;172;172mv7rrrrr7L..\033[38;2;252;238;238mB                    ");
// $display("\033[38;2;252;238;238m                                                        .::7L7rriiiirr77rrrrrrrr72BBBBBBBBBBBBvi:..  \033[38;2;252;172;172m.  \033[38;2;252;238;238mBr \033[38;2;252;172;172m77rrrrrvi \033[38;2;252;238;238mKi                    ");
// $display("\033[38;2;252;238;238m                                                    :rv7i::...........    .:i7BBBBQbPPPqPPPdEZQBBBBBr:.\033[38;2;252;238;238m ii \033[38;2;252;172;172mvvrrrrvr \033[38;2;252;238;238mvs                     ");
// $display("\033[38;2;252;238;238m                    .S77L.                      .rvi:. ..:r7QBBBBBBBBBBBgri.    .:BBBPqqKKqqqqPPPPPEQBBBZi  \033[38;2;252;172;172m:777vi \033[38;2;252;238;238mvI                      ");
// $display("\033[38;2;252;238;238m                    B: ..Jv                   isi. .:rBBBBBQZPPPPqqqPPdERBBBBBi.    :BBRKqqqqqqqqqqqqPKDDBB:  \033[38;2;252;172;172m:7. \033[38;2;252;238;238mJr                       ");
// $display("\033[38;2;252;238;238m                   vv SB: iu                rL: .iBBBQEPqqPPqqqqqqqqqqqqqPPPPbQBBB:   .EBQKqqqqqqPPPqqKqPPgBB:  .B:                        ");
// $display("\033[38;2;252;238;238m                  :R  BgBL..s7            rU: .qBBEKPqqqqqqqqqqqqqqqqqqqqqqqqqPPPEBBB:   EBEPPPEgQBBQEPqqqqKEBB: .s                        ");
// $display("\033[38;2;252;238;238m               .U7.  iBZBBBi :ji         5r .MBQqPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPKgBB:  .BBBBBdJrrSBBQKqqqqKZB7  I:                      ");
// $display("\033[38;2;252;238;238m              v2. :rBBBB: .BB:.ru7:    :5. rBQqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPPBB:  :.        .5BKqqqqqqBB. Kr                     ");
// $display("\033[38;2;252;238;238m             .B .BBQBB.   .RBBr  :L77ri2  BBqPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPbBB   \033[38;2;252;172;172m.irrrrri  \033[38;2;252;238;238mQQqqqqqqKRB. 2i                    ");
// $display("\033[38;2;252;238;238m              27 :BBU  rBBBdB \033[38;2;252;172;172m iri::::: \033[38;2;252;238;238m.BQKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqKRBs\033[38;2;252;172;172mirrr7777L: \033[38;2;252;238;238m7BqqqqqqqXZB. BLv772i              ");
// $display("\033[38;2;252;238;238m               rY  PK  .:dPMB \033[38;2;252;172;172m.Y77777r.\033[38;2;252;238;238m:BEqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPPBqi\033[38;2;252;172;172mirrrrrv: \033[38;2;252;238;238muBqqqqqqqqqgB  :.:. B:             ");
// $display("\033[38;2;252;238;238m                iu 7BBi  rMgB \033[38;2;252;172;172m.vrrrrri\033[38;2;252;238;238mrBEqKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQgi\033[38;2;252;172;172mirrrrv. \033[38;2;252;238;238mQQqqqqqqqqqXBb .BBB .s:.           ");
// $display("\033[38;2;252;238;238m                i7 BBdBBBPqbB \033[38;2;252;172;172m.vrrrri\033[38;2;252;238;238miDgPPbPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQDi\033[38;2;252;172;172mirr77 \033[38;2;252;238;238m:BdqqqqqqqqqqPB. rBB. .:iu7         ");
// $display("\033[38;2;252;238;238m                iX.:iBRKPqKXB.\033[38;2;252;172;172m 77rrr\033[38;2;252;238;238mi7QPBBBBPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPB7i\033[38;2;252;172;172mrr7r \033[38;2;252;238;238m.vBBPPqqqqqqKqBZ  BPBgri: 1B        ");
// $display("\033[38;2;252;238;238m                 ivr .BBqqKXBi \033[38;2;252;172;172mr7rri\033[38;2;252;238;238miQgQi   QZKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPEQi\033[38;2;252;172;172mirr7r.  \033[38;2;252;238;238miBBqPqqqqqqPB:.QPPRBBB LK        ");
// $display("\033[38;2;252;238;238m                   :I. iBgqgBZ \033[38;2;252;172;172m:7rr\033[38;2;252;238;238miJQPB.   gRqqqqqqqqPPPPPPPPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQ7\033[38;2;252;172;172mirrr7vr.  \033[38;2;252;238;238mUBqqPPgBBQPBBKqqqKB  B         ");
// $display("\033[38;2;252;238;238m                     v7 .BBR: \033[38;2;252;172;172m.r7ri\033[38;2;252;238;238miggqPBrrBBBBBBBBBBBBBBBBBBQEPPqqPPPqqqqqqqqqqqqqqqqqqqqqqqqqPgPi\033[38;2;252;172;172mirrrr7v7  \033[38;2;252;238;238mrBPBBP:.LBbPqqqqqB. u.        ");
// $display("\033[38;2;252;238;238m                      .j. . \033[38;2;252;172;172m :77rr\033[38;2;252;238;238miiBPqPbBB::::::.....:::iirrSBBBBBBBQZPPPPPqqqqqqqqqqqqqqqqqqqqEQi\033[38;2;252;172;172mirrrrrr7v \033[38;2;252;238;238m.BB:     :BPqqqqqDB .B        ");
// $display("\033[38;2;252;238;238m                       YL \033[38;2;252;172;172m.i77rrrr\033[38;2;252;238;238miLQPqqKQJ. \033[38;2;252;172;172m ............       \033[38;2;252;238;238m..:irBBBBBBZPPPqqqqqqqPPBBEPqqqdRr\033[38;2;252;172;172mirrrrrr7v \033[38;2;252;238;238m.B  .iBB  dQPqqqqPBi Y:       ");
// $display("\033[38;2;252;238;238m                     :U:.\033[38;2;252;172;172mrv7rrrrri\033[38;2;252;238;238miPgqqqqKZB.\033[38;2;252;172;172m.v77777777777777ri::..   \033[38;2;252;238;238m  ..:rBBBBQPPqqqqPBUvBEqqqPRr\033[38;2;252;172;172mirrrrrrvi\033[38;2;252;238;238m iB:RBBbB7 :BQqPqKqBR r7       ");
// $display("\033[38;2;252;238;238m                    iI.\033[38;2;252;172;172m.v7rrrrrrri\033[38;2;252;238;238midgqqqqqKB:\033[38;2;252;172;172m 77rrrrrrrrrrrrr77777777ri:..   \033[38;2;252;238;238m .:1BBBEPPB:   BbqqPQr\033[38;2;252;172;172mirrrr7vr\033[38;2;252;238;238m .BBBZPqqDB  .JBbqKPBi vi       ");
// $display("\033[38;2;252;238;238m                   :B \033[38;2;252;172;172miL7rrrrrrrri\033[38;2;252;238;238mibgqqqqqqBr\033[38;2;252;172;172m r7rrrrrrrrrrrrrrrrrrrrr777777ri:.  \033[38;2;252;238;238m .iBBBBi  .BbqqdRr\033[38;2;252;172;172mirr7v7: \033[38;2;252;238;238m.Bi.dBBPqqgB:  :BPqgB  B        ");
// $display("\033[38;2;252;238;238m                   .K.i\033[38;2;252;172;172mv7rrrrrrrri\033[38;2;252;238;238miZgqqqqqqEB \033[38;2;252;172;172m.vrrrrrrrrrrrrrrrrrrrrrrrrrrr777vv7i.  \033[38;2;252;238;238m :PBBBBPqqqEQ\033[38;2;252;172;172miir77:  \033[38;2;252;238;238m:BB:  .rBPqqEBB. iBZB. Rr        ");
// $display("\033[38;2;252;238;238m                    iM.:\033[38;2;252;172;172mv7rrrrrrrri\033[38;2;252;238;238mUQPqqqqqPBi\033[38;2;252;172;172m i7rrrrrrrrrrrrrrrrrrrrrrrrr77777i.   \033[38;2;252;238;238m.  :BddPqqqqEg\033[38;2;252;172;172miir7. \033[38;2;252;238;238mrBBPqBBP. :BXKqgB  BBB. 2r         ");
// $display("\033[38;2;252;238;238m                     :U:.\033[38;2;252;172;172miv77rrrrri\033[38;2;252;238;238mrBPqqqqqqPB: \033[38;2;252;172;172m:7777rrrrrrrrrrrrrrr777777ri.   \033[38;2;252;238;238m.:uBBBBZPqqqqqqPQL\033[38;2;252;172;172mirr77 \033[38;2;252;238;238m.BZqqPB:  qMqqPB. Yv:  Ur          ");
// $display("\033[38;2;252;238;238m                       1L:.\033[38;2;252;172;172m:77v77rii\033[38;2;252;238;238mqQPqqqqqPbBi \033[38;2;252;172;172m .ir777777777777777ri:..   \033[38;2;252;238;238m.:rBBBRPPPPPqqqqqqqgQ\033[38;2;252;172;172miirr7vr \033[38;2;252;238;238m:BqXQ: .BQPZBBq ...:vv.           ");
// $display("\033[38;2;252;238;238m                         LJi..\033[38;2;252;172;172m::r7rii\033[38;2;252;238;238mRgKPPPPqPqBB:.  \033[38;2;252;172;172m ............     \033[38;2;252;238;238m..:rBBBBPPqqKKKKqqqPPqPbB1\033[38;2;252;172;172mrvvvvvr  \033[38;2;252;238;238mBEEDQBBBBBRri. 7JLi              ");
// $display("\033[38;2;252;238;238m                           .jL\033[38;2;252;172;172m  777rrr\033[38;2;252;238;238mBBBBBBgEPPEBBBvri:::::::::irrrbBBBBBBDPPPPqqqqqqXPPZQBBBBr\033[38;2;252;172;172m.......\033[38;2;252;238;238m.:BBBBg1ri:....:rIr                 ");
// $display("\033[38;2;252;238;238m                            vI \033[38;2;252;172;172m:irrr:....\033[38;2;252;238;238m:rrEBBBBBBBBBBBBBBBBBBBBBBBBBBBBBQQBBBBBBBBBBBBBQr\033[38;2;252;172;172mi:...:.   \033[38;2;252;238;238m.:ii:.. .:.:irri::                    ");
// $display("\033[38;2;252;238;238m                             71vi\033[38;2;252;172;172m:::irrr::....\033[38;2;252;238;238m    ...:..::::irrr7777777777777rrii::....  ..::irvrr7sUJYv7777v7ii..                         ");
// $display("\033[38;2;252;238;238m                               .i777i. ..:rrri77rriiiiiii:::::::...............:::iiirr7vrrr:.                                             ");
// $display("\033[38;2;252;238;238m                                                      .::::::::::::::::::::::::::::::                                                      \033[m");
end endtask

task JohnCena; begin
$display("\033[48;2;100;100;103m \033[48;2;106;106;108m \033[48;2;100;100;105m \033[48;2;102;100;105m \033[48;2;106;103;108m \033[48;2;107;102;108m \033[48;2;108;103;109m \033[48;2;113;108;114m \033[48;2;116;111;117m \033[48;2;117;112;118m \033[48;2;118;113;119m \033[48;2;117;115;120m \033[48;2;118;116;121m \033[48;2;122;120;125m \033[48;2;125;123;128m \033[48;2;124;122;127m \033[48;2;124;122;127m \033[48;2;126;123;128m \033[48;2;125;123;127m \033[48;2;124;123;128m \033[48;2;119;122;129m \033[48;2;113;116;123m \033[48;2;97;100;107m \033[48;2;90;94;100m \033[48;2;88;93;99m \033[48;2;85;90;96m \033[48;2;80;85;91m \033[48;2;82;87;93m \033[48;2;80;85;91m \033[48;2;74;79;85m \033[48;2;70;75;80m \033[48;2;68;73;79m \033[48;2;67;72;78m \033[48;2;67;72;76m \033[48;2;66;71;77m \033[48;2;66;70;78m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;66;70;79m \033[48;2;65;69;78m \033[48;2;66;70;79m \033[48;2;68;72;83m \033[48;2;68;72;83m \033[48;2;66;70;81m \033[48;2;63;67;78m \033[48;2;60;64;75m \033[48;2;60;64;75m \033[48;2;59;63;74m \033[48;2;59;63;74m \033[48;2;59;63;74m \033[48;2;60;64;75m \033[48;2;60;64;75m \033[48;2;63;67;78m \033[48;2;65;69;80m \033[48;2;67;71;82m \033[48;2;69;73;82m \033[48;2;68;72;81m \033[48;2;68;72;83m \033[48;2;68;72;83m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;66;70;81m \033[48;2;67;71;82m \033[48;2;67;71;82m \033[48;2;65;72;82m \033[48;2;67;71;82m \033[48;2;68;72;83m \033[48;2;70;72;84m \033[48;2;73;74;86m \033[48;2;75;75;85m \033[48;2;76;76;86m \033[48;2;76;76;86m \033[48;2;76;76;86m \033[48;2;76;76;86m \033[48;2;76;76;86m \033[48;2;74;77;86m \033[48;2;74;77;86m \033[48;2;74;77;86m \033[48;2;73;77;86m \033[48;2;74;77;86m \033[48;2;77;78;87m \033[48;2;76;76;86m \033[48;2;77;74;85m \033[48;2;76;73;82m \033[48;2;76;73;82m \033[48;2;77;74;80m \033[48;2;78;74;81m \033[48;2;80;75;81m \033[48;2;79;74;80m \033[48;2;79;74;80m \033[48;2;79;74;80m \033[48;2;77;72;78m \033[48;2;76;71;77m \033[48;2;76;71;77m \033[48;2;76;71;77m \033[48;2;75;71;77m \033[48;2;73;70;77m \033[48;2;72;69;76m \033[48;2;69;66;73m \033[48;2;67;64;71m \033[48;2;69;64;71m \033[48;2;68;63;70m \033[48;2;66;61;68m \033[48;2;66;61;68m \033[48;2;64;61;66m \033[m");
$display("\033[48;2;112;110;115m \033[48;2;115;113;118m \033[48;2;115;113;118m \033[48;2;114;112;117m \033[48;2;116;114;119m \033[48;2;116;114;119m \033[48;2;117;112;118m \033[48;2;117;112;118m \033[48;2;119;115;120m \033[48;2;124;119;125m \033[48;2;129;124;130m \033[48;2;130;125;131m \033[48;2;131;126;132m \033[48;2;135;130;136m \033[48;2;142;137;143m \033[48;2;145;143;148m \033[48;2;145;143;148m \033[48;2;142;140;145m \033[48;2;142;140;145m \033[48;2;136;135;140m \033[48;2;131;131;139m \033[48;2;113;116;123m \033[48;2;98;101;108m \033[48;2;90;95;101m \033[48;2;88;91;98m \033[48;2;86;89;96m \033[48;2;83;87;94m \033[48;2;81;86;92m \033[48;2;74;79;85m \033[48;2;72;75;82m \033[48;2;69;72;79m \033[48;2;68;71;78m \033[48;2;67;70;77m \033[48;2;66;69;76m \033[48;2;66;69;76m \033[48;2;65;68;77m \033[48;2;64;67;76m \033[48;2;64;67;76m \033[48;2;64;68;77m \033[48;2;64;68;77m \033[48;2;66;70;79m \033[48;2;67;71;80m \033[48;2;64;68;77m \033[48;2;55;59;67m \033[48;2;50;54;63m \033[48;2;50;54;63m \033[48;2;50;54;63m \033[48;2;46;50;59m \033[48;2;46;50;59m \033[48;2;45;49;60m \033[48;2;45;49;60m \033[48;2;46;50;59m \033[48;2;47;51;60m \033[48;2;48;52;61m \033[48;2;48;52;62m \033[48;2;49;53;63m \033[48;2;53;57;68m \033[48;2;54;58;68m \033[48;2;52;56;67m \033[48;2;54;58;69m \033[48;2;64;68;79m \033[48;2;66;70;81m \033[48;2;65;69;80m \033[48;2;66;70;81m \033[48;2;67;70;82m \033[48;2;66;68;80m \033[48;2;66;68;80m \033[48;2;66;68;80m \033[48;2;66;68;80m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;65;69;79m \033[48;2;68;71;78m \033[48;2;69;72;79m \033[48;2;70;73;80m \033[48;2;71;74;81m \033[48;2;69;73;82m \033[48;2;69;73;82m \033[48;2;71;75;84m \033[48;2;69;76;84m \033[48;2;71;75;84m \033[48;2;70;73;82m \033[48;2;70;73;82m \033[48;2;72;72;83m \033[48;2;72;72;82m \033[48;2;72;70;81m \033[48;2;72;70;81m \033[48;2;72;69;78m \033[48;2;72;69;78m \033[48;2;74;68;77m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;75;70;77m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;74;69;76m \033[48;2;73;70;77m \033[48;2;72;69;76m \033[48;2;67;64;71m \033[48;2;66;63;70m \033[48;2;65;62;69m \033[48;2;64;61;68m \033[48;2;62;57;64m \033[48;2;60;54;62m \033[48;2;57;53;59m \033[m");
$display("\033[48;2;110;108;109m \033[48;2;112;111;111m \033[48;2;116;114;117m \033[48;2;124;122;125m \033[48;2;129;127;130m \033[48;2;129;127;130m \033[48;2;130;128;131m \033[48;2;130;128;131m \033[48;2;128;126;129m \033[48;2;128;126;129m \033[48;2;129;127;130m \033[48;2;131;129;134m \033[48;2;137;135;140m \033[48;2;139;137;142m \033[48;2;140;138;143m \033[48;2;142;142;146m \033[48;2;147;146;151m \033[48;2;144;144;148m \033[48;2;139;138;143m \033[48;2;130;130;135m \033[48;2;120;121;126m \033[48;2;98;102;107m \033[48;2;94;97;101m \033[48;2;86;91;95m \033[48;2;85;88;95m \033[48;2;83;86;93m \033[48;2;79;84;90m \033[48;2;77;82;88m \033[48;2;71;76;82m \033[48;2;70;75;81m \033[48;2;67;72;78m \033[48;2;66;71;77m \033[48;2;64;69;75m \033[48;2;64;69;73m \033[48;2;64;69;75m \033[48;2;65;69;77m \033[48;2;64;68;78m \033[48;2;64;68;77m \033[48;2;65;69;78m \033[48;2;65;69;78m \033[48;2;62;66;74m \033[48;2;53;57;66m \033[48;2;51;55;64m \033[48;2;50;54;63m \033[48;2;43;47;56m \033[48;2;43;47;56m \033[48;2;45;48;57m \033[48;2;43;48;55m \033[48;2;43;47;56m \033[48;2;44;48;57m \033[48;2;44;48;59m \033[48;2;44;47;59m \033[48;2;45;48;60m \033[48;2;47;50;62m \033[48;2;47;51;62m \033[48;2;48;51;63m \033[48;2;47;51;62m \033[48;2;48;51;62m \033[48;2;48;52;63m \033[48;2;46;50;61m \033[48;2;48;51;62m \033[48;2;50;54;65m \033[48;2;49;52;63m \033[48;2;53;57;68m \033[48;2;59;63;73m \033[48;2;63;68;79m \033[48;2;64;68;79m \033[48;2;65;69;80m \033[48;2;65;69;80m \033[48;2;64;68;78m \033[48;2;64;68;78m \033[48;2;64;68;78m \033[48;2;64;68;78m \033[48;2;64;69;78m \033[48;2;64;69;75m \033[48;2;65;70;76m \033[48;2;65;70;76m \033[48;2;67;72;78m \033[48;2;67;72;80m \033[48;2;67;72;80m \033[48;2;68;72;80m \033[48;2;69;72;80m \033[48;2;69;72;81m \033[48;2;70;72;81m \033[48;2;72;72;81m \033[48;2;72;70;80m \033[48;2;70;69;79m \033[48;2;70;68;79m \033[48;2;69;67;78m \033[48;2;71;68;78m \033[48;2;72;68;78m \033[48;2;72;68;75m \033[48;2;70;67;74m \033[48;2;70;67;74m \033[48;2;71;68;75m \033[48;2;71;68;75m \033[48;2;69;67;73m \033[48;2;68;65;72m \033[48;2;67;64;72m \033[48;2;67;64;72m \033[48;2;68;64;72m \033[48;2;68;63;70m \033[48;2;68;63;70m \033[48;2;67;62;69m \033[48;2;67;61;68m \033[48;2;64;62;67m \033[48;2;64;59;65m \033[48;2;61;56;62m \033[48;2;60;53;60m \033[48;2;58;51;58m \033[m");
$display("\033[48;2;96;95;91m \033[48;2;98;97;93m \033[48;2;104;102;103m \033[48;2;104;102;103m \033[48;2;109;107;108m \033[48;2;109;107;108m \033[48;2;112;113;112m \033[48;2;116;116;116m \033[48;2;117;117;117m \033[48;2;119;120;119m \033[48;2;122;122;124m \033[48;2;120;119;124m \033[48;2;121;120;125m \033[48;2;119;118;123m \033[48;2;123;121;127m \033[48;2;124;128;130m \033[48;2;124;128;131m \033[48;2;130;134;137m \033[48;2;123;127;130m \033[48;2;116;121;125m \033[48;2;101;102;106m \033[48;2;89;94;96m \033[48;2;85;89;92m \033[48;2;82;87;90m \033[48;2;82;85;92m \033[48;2;80;83;90m \033[48;2;73;77;84m \033[48;2;70;75;81m \033[48;2;68;73;79m \033[48;2;68;71;78m \033[48;2;66;69;76m \033[48;2;65;68;75m \033[48;2;64;67;74m \033[48;2;63;66;73m \033[48;2;64;67;74m \033[48;2;64;68;77m \033[48;2;65;68;77m \033[48;2;65;68;77m \033[48;2;66;68;78m \033[48;2;59;61;70m \033[48;2;50;52;61m \033[48;2;44;46;55m \033[48;2;43;46;55m \033[48;2;41;44;53m \033[48;2;44;46;55m \033[48;2;43;46;54m \033[48;2;43;45;54m \033[48;2;43;45;54m \033[48;2;43;46;56m \033[48;2;42;44;54m \033[48;2;43;45;57m \033[48;2;45;47;60m \033[48;2;46;48;61m \033[48;2;46;48;61m \033[48;2;46;48;61m \033[48;2;47;49;62m \033[48;2;48;49;61m \033[48;2;46;48;60m \033[48;2;46;47;59m \033[48;2;45;47;59m \033[48;2;48;49;61m \033[48;2;46;48;60m \033[48;2;45;48;59m \033[48;2;45;47;59m \033[48;2;46;48;60m \033[48;2;53;55;67m \033[48;2;54;56;68m \033[48;2;62;64;76m \033[48;2;62;64;76m \033[48;2;62;65;74m \033[48;2;61;65;74m \033[48;2;61;65;74m \033[48;2;61;65;74m \033[48;2;61;65;74m \033[48;2;63;67;74m \033[48;2;63;66;74m \033[48;2;65;68;75m \033[48;2;65;67;75m \033[48;2;63;68;74m \033[48;2;64;69;75m \033[48;2;67;67;75m \033[48;2;69;67;75m \033[48;2;68;68;76m \033[48;2;69;68;76m \033[48;2;69;68;76m \033[48;2;70;67;76m \033[48;2;69;66;75m \033[48;2;68;66;77m \033[48;2;68;66;77m \033[48;2;68;65;74m \033[48;2;68;65;74m \033[48;2;67;64;73m \033[48;2;66;65;71m \033[48;2;66;65;71m \033[48;2;65;63;70m \033[48;2;65;63;70m \033[48;2;65;64;70m \033[48;2;64;63;69m \033[48;2;64;62;68m \033[48;2;63;62;68m \033[48;2;65;61;68m \033[48;2;67;60;67m \033[48;2;66;59;67m \033[48;2;66;59;67m \033[48;2;66;59;67m \033[48;2;64;57;65m \033[48;2;62;55;63m \033[48;2;63;52;62m \033[48;2;61;51;61m \033[48;2;58;51;58m \033[m");
$display("\033[48;2;66;66;66m \033[48;2;66;65;66m \033[48;2;73;71;74m \033[48;2;78;76;79m \033[48;2;81;79;82m \033[48;2;86;84;87m \033[48;2;86;86;88m \033[48;2;87;87;89m \033[48;2;90;90;92m \033[48;2;95;95;97m \033[48;2;99;99;101m \033[48;2;100;101;103m \033[48;2;102;104;106m \033[48;2;105;107;109m \033[48;2;109;112;113m \033[48;2;114;118;119m \033[48;2;122;126;127m \033[48;2;129;133;134m \033[48;2;123;127;128m \033[48;2;114;118;119m \033[48;2;103;107;110m \033[48;2;93;97;100m \033[48;2;88;91;96m \033[48;2;87;90;95m \033[48;2;85;87;92m \033[48;2;81;83;88m \033[48;2;76;78;85m \033[48;2;74;75;83m \033[48;2;71;73;82m \033[48;2;70;70;78m \033[48;2;69;69;77m \033[48;2;68;67;75m \033[48;2;68;67;75m \033[48;2;68;68;78m \033[48;2;67;67;77m \033[48;2;86;86;96m \033[48;2;71;71;81m \033[48;2;51;51;61m \033[48;2;48;46;59m \033[48;2;46;44;57m \033[48;2;46;44;57m \033[48;2;43;41;54m \033[48;2;42;40;53m \033[48;2;43;41;54m \033[48;2;45;43;56m \033[48;2;45;43;56m \033[48;2;45;43;56m \033[48;2;47;43;57m \033[48;2;47;44;58m \033[48;2;47;45;58m \033[48;2;49;47;60m \033[48;2;49;49;61m \033[48;2;49;49;61m \033[48;2;49;47;60m \033[48;2;49;47;60m \033[48;2;50;46;60m \033[48;2;50;46;60m \033[48;2;50;46;60m \033[48;2;50;46;60m \033[48;2;50;46;60m \033[48;2;48;44;58m \033[48;2;48;44;58m \033[48;2;47;45;58m \033[48;2;47;45;58m \033[48;2;47;45;58m \033[48;2;43;41;54m \033[48;2;42;40;53m \033[48;2;46;44;55m \033[48;2;58;56;67m \033[48;2;60;61;71m \033[48;2;61;61;71m \033[48;2;61;61;71m \033[48;2;63;61;72m \033[48;2;63;61;72m \033[48;2;62;62;72m \033[48;2;62;62;72m \033[48;2;64;62;73m \033[48;2;64;62;73m \033[48;2;64;64;72m \033[48;2;64;64;72m \033[48;2;66;66;74m \033[48;2;65;65;73m \033[48;2;65;66;74m \033[48;2;66;65;73m \033[48;2;66;65;73m \033[48;2;67;66;74m \033[48;2;66;65;73m \033[48;2;65;63;74m \033[48;2;65;64;72m \033[48;2;65;62;71m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;62;59;66m \033[48;2;62;59;66m \033[48;2;63;59;66m \033[48;2;64;59;66m \033[48;2;64;59;66m \033[48;2;63;58;65m \033[48;2;62;57;64m \033[48;2;62;57;63m \033[48;2;60;55;61m \033[48;2;58;51;58m \033[48;2;57;50;57m \033[48;2;54;49;54m \033[m");
$display("\033[48;2;61;61;61m \033[48;2;58;59;59m \033[48;2;60;58;61m \033[48;2;60;58;61m \033[48;2;62;60;63m \033[48;2;65;63;66m \033[48;2;64;64;66m \033[48;2;72;72;74m \033[48;2;74;74;76m \033[48;2;79;79;81m \033[48;2;83;84;86m \033[48;2;85;91;91m \033[48;2;89;96;95m \033[48;2;93;100;99m \033[48;2;99;106;106m \033[48;2;106;112;112m \033[48;2;115;121;121m \033[48;2;123;129;129m \033[48;2;124;130;130m \033[48;2;126;132;132m \033[48;2;123;127;126m \033[48;2;114;118;119m \033[48;2;107;111;113m \033[48;2;100;104;107m \033[48;2;91;96;100m \033[48;2;83;88;91m \033[48;2;77;82;88m \033[48;2;74;79;85m \033[48;2;72;76;85m \033[48;2;71;71;81m \033[48;2;69;69;79m \033[48;2;69;67;78m \033[48;2;69;67;78m \033[48;2;69;67;78m \033[48;2;75;73;84m \033[48;2;62;60;71m \033[48;2;50;48;59m \033[48;2;46;44;55m \033[48;2;47;47;57m \033[48;2;46;46;56m \033[48;2;46;46;56m \033[48;2;47;47;57m \033[48;2;48;46;59m \033[48;2;49;47;60m \033[48;2;50;48;61m \033[48;2;50;48;61m \033[48;2;50;47;60m \033[48;2;50;44;59m \033[48;2;52;46;60m \033[48;2;52;48;62m \033[48;2;51;47;62m \033[48;2;52;50;63m \033[48;2;51;49;62m \033[48;2;51;47;61m \033[48;2;50;46;60m \033[48;2;52;46;60m \033[48;2;52;44;59m \033[48;2;52;44;59m \033[48;2;52;44;59m \033[48;2;51;43;58m \033[48;2;50;44;58m \033[48;2;48;42;56m \033[48;2;44;40;54m \033[48;2;44;40;54m \033[48;2;43;41;54m \033[48;2;44;40;54m \033[48;2;43;39;53m \033[48;2;44;41;52m \033[48;2;44;41;52m \033[48;2;48;45;56m \033[48;2;57;55;66m \033[48;2;57;58;67m \033[48;2;59;60;70m \033[48;2;60;63;72m \033[48;2;59;62;71m \033[48;2;59;62;71m \033[48;2;61;61;71m \033[48;2;62;62;72m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;64;63;71m \033[48;2;64;63;71m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;61;72m \033[48;2;63;62;70m \033[48;2;64;61;70m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;61;58;65m \033[48;2;60;57;64m \033[48;2;62;57;64m \033[48;2;61;56;63m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;59;54;60m \033[48;2;59;54;60m \033[48;2;59;54;60m \033[48;2;59;54;60m \033[48;2;59;54;60m \033[48;2;59;54;60m \033[48;2;59;52;59m \033[48;2;57;50;57m \033[48;2;54;49;55m \033[m");
$display("\033[48;2;56;56;58m \033[48;2;55;55;57m \033[48;2;56;56;58m \033[48;2;56;56;58m \033[48;2;55;55;57m \033[48;2;49;49;50m \033[48;2;43;43;45m \033[48;2;44;44;45m \033[48;2;44;44;45m \033[48;2;60;60;62m \033[48;2;79;79;81m \033[48;2;85;86;89m \033[48;2;86;90;93m \033[48;2;91;95;98m \033[48;2;97;102;103m \033[48;2;106;112;112m \033[48;2;117;123;123m \033[48;2;148;152;153m \033[48;2;158;162;163m \033[48;2;168;171;172m \033[48;2;168;168;168m \033[48;2;159;159;159m \033[48;2;144;144;144m \033[48;2;128;128;128m \033[48;2;106;109;113m \033[48;2;89;92;96m \033[48;2;82;87;93m \033[48;2;78;83;89m \033[48;2;75;79;87m \033[48;2;74;76;86m \033[48;2;73;73;83m \033[48;2;75;73;84m \033[48;2;76;74;85m \033[48;2;80;77;92m \033[48;2;70;68;80m \033[48;2;57;55;66m \033[48;2;51;50;59m \033[48;2;50;49;57m \033[48;2;48;48;56m \033[48;2;49;48;56m \033[48;2;52;50;60m \033[48;2;57;54;64m \033[48;2;59;56;63m \033[48;2;61;57;64m \033[48;2;63;57;65m \033[48;2;64;59;65m \033[48;2;67;59;67m \033[48;2;71;61;69m \033[48;2;72;61;70m \033[48;2;73;61;71m \033[48;2;79;68;77m \033[48;2;76;67;75m \033[48;2;69;61;69m \033[48;2;68;58;66m \033[48;2;66;57;66m \033[48;2;59;50;58m \033[48;2;55;47;59m \033[48;2;53;44;56m \033[48;2;54;44;56m \033[48;2;54;42;56m \033[48;2;54;46;61m \033[48;2;48;42;56m \033[48;2;44;40;52m \033[48;2;42;40;51m \033[48;2;42;40;52m \033[48;2;43;38;51m \033[48;2;42;37;50m \033[48;2;42;37;50m \033[48;2;43;38;51m \033[48;2;45;40;52m \033[48;2;47;44;55m \033[48;2;54;52;63m \033[48;2;61;59;70m \033[48;2;62;60;71m \033[48;2;62;60;71m \033[48;2;62;60;71m \033[48;2;61;59;70m \033[48;2;62;60;71m \033[48;2;62;61;69m \033[48;2;63;62;70m \033[48;2;64;63;71m \033[48;2;64;63;71m \033[48;2;64;63;71m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;59;56;63m \033[48;2;59;56;63m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;59;54;60m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;59;54;60m \033[48;2;60;53;60m \033[48;2;59;52;59m \033[48;2;57;50;57m \033[48;2;56;49;57m \033[48;2;54;49;55m \033[m");
$display("\033[48;2;44;44;46m \033[48;2;46;46;48m \033[48;2;52;51;56m \033[48;2;68;67;72m \033[48;2;74;73;77m \033[48;2;74;73;77m \033[48;2;74;73;77m \033[48;2;72;71;76m \033[48;2;65;64;69m \033[48;2;60;59;64m \033[48;2;55;55;59m \033[48;2;57;58;63m \033[48;2;65;68;73m \033[48;2;98;101;106m \033[48;2;140;145;149m \033[48;2;222;226;227m \033[48;2;250;254;255m \033[48;2;252;254;255m \033[48;2;253;254;255m \033[48;2;252;253;255m \033[48;2;253;253;253m \033[48;2;255;255;255m \033[48;2;226;226;226m \033[48;2;160;160;160m \033[48;2;129;131;136m \033[48;2;106;109;115m \033[48;2;93;98;104m \033[48;2;88;92;99m \033[48;2;81;85;94m \033[48;2;78;80;88m \033[48;2;74;77;84m \033[48;2;76;77;85m \033[48;2;86;86;94m \033[48;2;74;72;83m \033[48;2;54;53;60m \033[48;2;45;44;52m \033[48;2;43;42;48m \033[48;2;40;39;45m \033[48;2;48;45;55m \033[48;2;60;55;62m \033[48;2;69;61;66m \033[48;2;74;63;67m \033[48;2;79;64;68m \033[48;2;82;66;69m \033[48;2;84;65;67m \033[48;2;90;66;70m \033[48;2;95;68;71m \033[48;2;101;70;75m \033[48;2;105;73;79m \033[48;2;109;78;83m \033[48;2;112;81;86m \033[48;2;113;82;86m \033[48;2;112;81;86m \033[48;2;110;80;85m \033[48;2;110;80;84m \033[48;2;109;79;83m \033[48;2;106;78;85m \033[48;2;102;76;82m \033[48;2;102;76;82m \033[48;2;97;73;78m \033[48;2;82;61;68m \033[48;2;69;51;58m \033[48;2;60;46;54m \033[48;2;52;43;51m \033[48;2;49;42;50m \033[48;2;46;40;47m \033[48;2;44;37;45m \033[48;2;44;37;45m \033[48;2;45;38;46m \033[48;2;45;37;50m \033[48;2;45;39;51m \033[48;2;46;40;52m \033[48;2;43;41;52m \033[48;2;57;54;65m \033[48;2;60;58;69m \033[48;2;61;59;70m \033[48;2;62;60;71m \033[48;2;63;61;72m \033[48;2;62;61;69m \033[48;2;62;61;69m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;62;70m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;61;57;65m \033[48;2;60;57;64m \033[48;2;60;57;64m \033[48;2;61;56;62m \033[48;2;60;55;61m \033[48;2;61;56;62m \033[48;2;61;56;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;61m \033[48;2;59;54;60m \033[48;2;58;53;59m \033[48;2;59;54;60m \033[48;2;58;53;59m \033[48;2;59;53;57m \033[48;2;59;53;57m \033[48;2;57;51;55m \033[48;2;56;50;54m \033[48;2;55;50;54m \033[m");
$display("\033[48;2;93;90;97m \033[48;2;93;90;98m \033[48;2;87;84;91m \033[48;2;87;84;91m \033[48;2;83;80;87m \033[48;2;79;76;83m \033[48;2;77;73;80m \033[48;2;76;73;80m \033[48;2;78;75;82m \033[48;2;75;72;79m \033[48;2;69;68;74m \033[48;2;59;62;67m \033[48;2;58;61;67m \033[48;2;65;68;73m \033[48;2;112;115;120m \033[48;2;207;212;212m \033[48;2;252;255;255m \033[48;2;253;255;254m \033[48;2;254;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;234;234;234m \033[48;2;155;161;161m \033[48;2;118;123;125m \033[48;2;101;106;108m \033[48;2;86;91;95m \033[48;2;78;83;87m \033[48;2;72;77;81m \033[48;2;70;75;79m \033[48;2;69;74;78m \033[48;2;56;61;65m \033[48;2;49;49;59m \033[48;2;41;41;49m \033[48;2;39;38;44m \033[48;2;37;36;41m \033[48;2;46;45;49m \033[48;2;69;61;66m \033[48;2;76;64;68m \033[48;2;81;63;66m \033[48;2;83;63;64m \033[48;2;85;62;60m \033[48;2;92;65;65m \033[48;2;103;72;70m \033[48;2;109;74;72m \033[48;2;115;76;75m \033[48;2;118;81;75m \033[48;2;125;85;80m \033[48;2;129;89;84m \033[48;2;133;92;87m \033[48;2;133;91;90m \033[48;2;133;91;90m \033[48;2;133;92;90m \033[48;2;133;91;90m \033[48;2;132;92;90m \033[48;2;136;91;93m \033[48;2;131;87;87m \033[48;2;127;85;86m \033[48;2;124;83;84m \033[48;2;115;79;79m \033[48;2;110;79;77m \033[48;2;105;75;77m \033[48;2;95;72;73m \033[48;2;81;61;63m \033[48;2;65;52;55m \033[48;2;48;39;43m \033[48;2;43;38;41m \033[48;2;43;38;42m \033[48;2;45;37;47m \033[48;2;45;39;49m \033[48;2;46;40;52m \033[48;2;41;38;49m \033[48;2;50;47;58m \033[48;2;62;60;71m \033[48;2;61;59;70m \033[48;2;63;61;72m \033[48;2;63;61;72m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;62;59;66m \033[48;2;61;58;65m \033[48;2;61;58;65m \033[48;2;60;57;64m \033[48;2;60;57;64m \033[48;2;61;57;64m \033[48;2;63;58;64m \033[48;2;62;57;63m \033[48;2;61;56;62m \033[48;2;61;56;62m \033[48;2;60;55;62m \033[48;2;60;55;61m \033[48;2;60;55;61m \033[48;2;60;55;59m \033[48;2;60;55;59m \033[48;2;60;54;58m \033[48;2;60;54;58m \033[48;2;60;54;58m \033[48;2;59;53;57m \033[48;2;58;53;59m \033[48;2;58;53;57m \033[48;2;56;51;55m \033[48;2;55;51;52m \033[48;2;55;51;52m \033[m");
$display("\033[48;2;59;57;63m \033[48;2;51;48;57m \033[48;2;39;36;44m \033[48;2;48;46;52m \033[48;2;60;57;64m \033[48;2;74;71;78m \033[48;2;76;75;81m \033[48;2;85;84;90m \033[48;2;79;78;83m \033[48;2;75;74;80m \033[48;2;76;75;81m \033[48;2;75;76;81m \033[48;2;75;76;81m \033[48;2;73;74;79m \033[48;2;80;81;86m \033[48;2;92;92;96m \033[48;2;150;151;155m \033[48;2;226;226;228m \033[48;2;254;254;255m \033[48;2;255;255;255m \033[48;2;255;254;252m \033[48;2;255;255;253m \033[48;2;253;252;250m \033[48;2;250;249;247m \033[48;2;154;158;161m \033[48;2;118;120;124m \033[48;2;95;97;102m \033[48;2;88;90;96m \033[48;2;83;83;91m \033[48;2;77;78;83m \033[48;2;72;73;78m \033[48;2;79;80;84m \033[48;2;71;72;77m \033[48;2;46;44;53m \033[48;2;38;35;42m \033[48;2;37;33;39m \033[48;2;40;35;39m \033[48;2;65;59;62m \033[48;2;79;64;67m \033[48;2;86;68;68m \033[48;2;90;67;65m \033[48;2;93;68;64m \033[48;2;102;73;65m \033[48;2;109;79;71m \033[48;2;121;85;77m \033[48;2;127;87;81m \033[48;2;134;91;84m \033[48;2;138;95;85m \033[48;2;145;98;90m \033[48;2;148;102;93m \033[48;2;153;104;97m \033[48;2;153;104;97m \033[48;2;154;105;99m \033[48;2;156;107;102m \033[48;2;153;104;98m \033[48;2;157;108;100m \033[48;2;157;107;98m \033[48;2;155;106;97m \033[48;2;155;107;97m \033[48;2;152;105;95m \033[48;2;143;98;93m \033[48;2;133;89;86m \033[48;2;125;85;83m \033[48;2;117;82;80m \033[48;2;107;77;75m \033[48;2;94;69;70m \033[48;2;79;63;64m \033[48;2;49;38;41m \033[48;2;48;39;44m \033[48;2;45;38;46m \033[48;2;44;39;46m \033[48;2;43;37;47m \033[48;2;39;36;45m \033[48;2;37;34;43m \033[48;2;56;53;62m \033[48;2;64;61;70m \033[48;2;64;61;70m \033[48;2;64;61;70m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;64;61;68m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;60;58;63m \033[48;2;60;58;63m \033[48;2;60;58;63m \033[48;2;60;58;63m \033[48;2;61;58;63m \033[48;2;63;58;64m \033[48;2;61;56;62m \033[48;2;61;56;62m \033[48;2;61;56;62m \033[48;2;60;55;62m \033[48;2;60;55;61m \033[48;2;59;54;60m \033[48;2;59;54;58m \033[48;2;59;54;58m \033[48;2;58;53;57m \033[48;2;58;53;57m \033[48;2;58;53;57m \033[48;2;58;53;57m \033[48;2;58;53;57m \033[48;2;58;54;55m \033[48;2;57;53;54m \033[48;2;56;52;51m \033[48;2;55;51;52m \033[m");
$display("\033[48;2;31;30;35m \033[48;2;32;29;36m \033[48;2;33;30;37m \033[48;2;42;39;45m \033[48;2;55;54;60m \033[48;2;73;72;78m \033[48;2;90;89;95m \033[48;2;90;89;95m \033[48;2;88;87;93m \033[48;2;59;58;65m \033[48;2;59;58;64m \033[48;2;70;69;75m \033[48;2;70;69;75m \033[48;2;73;72;78m \033[48;2;70;69;75m \033[48;2;82;81;87m \033[48;2;101;100;105m \033[48;2;141;141;144m \033[48;2;145;145;147m \033[48;2;147;146;146m \033[48;2;152;147;147m \033[48;2;152;148;145m \033[48;2;151;146;144m \033[48;2;141;137;132m \033[48;2;122;121;117m \033[48;2;109;104;102m \033[48;2;97;93;92m \033[48;2;94;88;88m \033[48;2;108;105;106m \033[48;2;77;75;76m \033[48;2;75;73;76m \033[48;2;86;84;89m \033[48;2;57;55;60m \033[48;2;47;40;50m \033[48;2;45;40;47m \033[48;2;44;39;40m \033[48;2;63;53;51m \033[48;2;82;68;67m \033[48;2;88;68;67m \033[48;2;96;71;69m \033[48;2;106;78;71m \033[48;2;113;83;74m \033[48;2;123;88;77m \033[48;2;126;90;78m \033[48;2;133;93;81m \033[48;2;140;96;82m \033[48;2;147;99;86m \033[48;2;154;102;91m \033[48;2;159;107;94m \033[48;2;164;110;99m \033[48;2;168;114;101m \033[48;2;181;127;115m \033[48;2;185;131;119m \033[48;2;191;137;124m \033[48;2;195;142;129m \033[48;2;192;138;127m \033[48;2;181;127;116m \033[48;2;178;124;114m \033[48;2;170;116;106m \033[48;2;166;113;101m \033[48;2;167;113;103m \033[48;2;161;109;101m \033[48;2;152;104;98m \033[48;2;141;96;92m \033[48;2;129;88;83m \033[48;2;118;81;78m \033[48;2;108;79;77m \033[48;2;86;64;67m \033[48;2;59;40;44m \033[48;2;47;34;41m \033[48;2;45;37;41m \033[48;2;41;39;44m \033[48;2;39;36;44m \033[48;2;40;34;44m \033[48;2;56;53;60m \033[48;2;63;59;67m \033[48;2;63;60;67m \033[48;2;62;59;66m \033[48;2;63;58;65m \033[48;2;63;58;65m \033[48;2;64;59;66m \033[48;2;64;59;66m \033[48;2;63;60;67m \033[48;2;61;58;65m \033[48;2;60;57;64m \033[48;2;61;57;63m \033[48;2;62;57;63m \033[48;2;62;57;63m \033[48;2;62;57;63m \033[48;2;61;56;62m \033[48;2;61;56;62m \033[48;2;60;55;61m \033[48;2;60;55;61m \033[48;2;59;54;60m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;56;51;57m \033[48;2;56;51;57m \033[48;2;54;52;57m \033[48;2;54;52;57m \033[48;2;54;52;57m \033[48;2;54;52;57m \033[48;2;54;52;57m \033[48;2;54;52;55m \033[48;2;54;52;55m \033[48;2;55;53;56m \033[48;2;55;53;53m \033[48;2;55;51;48m \033[48;2;56;51;48m \033[48;2;54;50;47m \033[m");
$display("\033[48;2;30;29;35m \033[48;2;30;29;34m \033[48;2;35;32;39m \033[48;2;67;64;71m \033[48;2;87;86;92m \033[48;2;90;89;95m \033[48;2;91;90;96m \033[48;2;91;90;96m \033[48;2;95;94;100m \033[48;2;95;94;100m \033[48;2;93;92;98m \033[48;2;94;93;98m \033[48;2;93;92;98m \033[48;2;90;89;96m \033[48;2;95;94;100m \033[48;2;101;100;106m \033[48;2;107;106;111m \033[48;2;121;121;121m \033[48;2;122;122;121m \033[48;2;123;123;121m \033[48;2;123;122;118m \033[48;2;124;123;118m \033[48;2;127;126;120m \033[48;2;126;126;118m \033[48;2;128;127;123m \033[48;2;131;130;126m \033[48;2;144;140;137m \033[48;2;149;145;142m \033[48;2;158;154;153m \033[48;2;154;153;151m \033[48;2;120;118;119m \033[48;2;86;84;88m \033[48;2;51;49;54m \033[48;2;46;38;49m \033[48;2;44;39;44m \033[48;2;58;49;50m \033[48;2;78;63;61m \033[48;2;93;75;70m \033[48;2;102;78;75m \033[48;2;113;86;79m \033[48;2;118;85;76m \033[48;2;124;90;78m \033[48;2;133;95;80m \033[48;2;136;96;80m \033[48;2;145;101;84m \033[48;2;151;104;88m \033[48;2;157;108;91m \033[48;2;166;113;99m \033[48;2;171;117;103m \033[48;2;177;121;106m \033[48;2;180;124;109m \033[48;2;181;124;107m \033[48;2;186;130;113m \033[48;2;190;134;117m \033[48;2;187;131;114m \033[48;2;192;135;118m \033[48;2;189;133;116m \033[48;2;182;127;111m \033[48;2;180;125;109m \033[48;2;177;121;104m \033[48;2;177;119;105m \033[48;2;172;116;103m \033[48;2;162;109;98m \033[48;2;153;103;95m \033[48;2;145;98;91m \033[48;2;130;89;81m \033[48;2;117;80;77m \033[48;2;100;70;70m \033[48;2;78;52;56m \033[48;2;52;33;39m \033[48;2;47;35;39m \033[48;2;42;37;43m \033[48;2;39;36;42m \033[48;2;37;34;41m \033[48;2;56;53;59m \033[48;2;63;60;66m \033[48;2;60;57;64m \033[48;2;59;56;63m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;60;55;62m \033[48;2;59;56;63m \033[48;2;57;56;62m \033[48;2;57;54;61m \033[48;2;57;53;59m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;58;53;59m \033[48;2;57;52;58m \033[48;2;57;52;58m \033[48;2;56;51;57m \033[48;2;55;50;56m \033[48;2;55;50;56m \033[48;2;53;48;54m \033[48;2;53;48;54m \033[48;2;51;49;54m \033[48;2;50;49;54m \033[48;2;50;49;54m \033[48;2;51;48;55m \033[48;2;51;49;54m \033[48;2;51;49;52m \033[48;2;51;49;52m \033[48;2;54;52;57m \033[48;2;53;51;51m \033[48;2;55;52;47m \033[48;2;56;51;48m \033[48;2;54;50;47m \033[m");
$display("\033[48;2;71;69;74m \033[48;2;78;76;82m \033[48;2;83;81;86m \033[48;2;93;91;96m \033[48;2;92;91;96m \033[48;2;93;92;97m \033[48;2;93;92;97m \033[48;2;94;93;98m \033[48;2;94;93;98m \033[48;2;95;94;99m \033[48;2;95;94;99m \033[48;2;95;94;99m \033[48;2;94;93;98m \033[48;2;95;94;99m \033[48;2;99;98;103m \033[48;2;103;104;105m \033[48;2;109;109;111m \033[48;2;116;116;114m \033[48;2;120;120;117m \033[48;2;135;136;131m \033[48;2;146;147;141m \033[48;2;158;159;151m \033[48;2;164;165;157m \033[48;2;157;159;148m \033[48;2;155;156;147m \033[48;2;159;160;152m \033[48;2;158;158;152m \033[48;2;169;168;163m \033[48;2;146;145;142m \033[48;2;138;137;134m \033[48;2;131;129;130m \033[48;2;79;78;82m \033[48;2;39;37;42m \033[48;2;45;38;46m \033[48;2;45;39;43m \033[48;2;73;61;61m \033[48;2;94;73;72m \033[48;2;104;79;74m \033[48;2;112;85;78m \033[48;2;119;89;79m \033[48;2;129;95;83m \033[48;2;136;98;84m \033[48;2;146;105;87m \033[48;2;150;108;91m \033[48;2;160;113;93m \033[48;2;166;116;96m \033[48;2;171;120;99m \033[48;2;183;128;110m \033[48;2;188;132;115m \033[48;2;189;132;113m \033[48;2;191;134;115m \033[48;2;193;135;113m \033[48;2;197;139;117m \033[48;2;200;142;120m \033[48;2;199;141;119m \033[48;2;193;135;112m \033[48;2;191;133;110m \033[48;2;192;134;110m \033[48;2;191;133;109m \033[48;2;188;130;106m \033[48;2;187;126;105m \033[48;2;179;121;101m \033[48;2;172;116;99m \033[48;2;164;111;96m \033[48;2;158;106;93m \033[48;2;147;99;87m \033[48;2;132;89;82m \033[48;2;120;84;79m \033[48;2;100;69;66m \033[48;2;57;33;39m \033[48;2;49;35;37m \033[48;2;40;35;39m \033[48;2;35;34;38m \033[48;2;35;34;39m \033[48;2;56;54;59m \033[48;2;60;58;63m \033[48;2;60;58;63m \033[48;2;58;56;61m \033[48;2;59;54;61m \033[48;2;59;54;61m \033[48;2;58;53;60m \033[48;2;57;52;59m \033[48;2;55;52;59m \033[48;2;53;50;57m \033[48;2;53;50;57m \033[48;2;53;49;54m \033[48;2;52;47;53m \033[48;2;52;47;53m \033[48;2;51;46;52m \033[48;2;51;46;52m \033[48;2;51;46;52m \033[48;2;51;46;52m \033[48;2;52;47;53m \033[48;2;52;47;53m \033[48;2;50;45;51m \033[48;2;50;45;51m \033[48;2;51;46;52m \033[48;2;51;46;52m \033[48;2;49;47;52m \033[48;2;49;47;52m \033[48;2;49;47;53m \033[48;2;50;47;54m \033[48;2;50;48;53m \033[48;2;50;48;51m \033[48;2;50;48;51m \033[48;2;50;48;53m \033[48;2;51;50;50m \033[48;2;54;52;47m \033[48;2;54;50;46m \033[48;2;52;49;46m \033[m");
$display("\033[48;2;83;81;84m \033[48;2;92;90;93m \033[48;2;94;90;96m \033[48;2;96;92;98m \033[48;2;96;93;97m \033[48;2;98;94;98m \033[48;2;98;96;99m \033[48;2;98;96;99m \033[48;2;98;96;99m \033[48;2;98;96;99m \033[48;2;97;95;98m \033[48;2;97;95;98m \033[48;2;98;96;99m \033[48;2;98;96;97m \033[48;2;101;99;100m \033[48;2;107;106;103m \033[48;2;112;111;108m \033[48;2;122;121;118m \033[48;2;132;131;129m \033[48;2;148;147;144m \033[48;2;147;145;146m \033[48;2;150;149;147m \033[48;2;156;155;150m \033[48;2;146;145;140m \033[48;2;134;135;130m \033[48;2;135;136;131m \033[48;2;126;125;121m \033[48;2;124;123;119m \033[48;2;122;121;117m \033[48;2;110;109;107m \033[48;2;107;103;108m \033[48;2;80;75;81m \033[48;2;42;35;41m \033[48;2;46;40;42m \033[48;2;73;61;63m \033[48;2;90;72;71m \033[48;2;97;73;67m \033[48;2;106;79;72m \033[48;2;112;83;74m \033[48;2;122;89;79m \033[48;2;134;98;86m \033[48;2;145;107;95m \033[48;2;153;111;95m \033[48;2;167;124;108m \033[48;2;174;129;110m \033[48;2;179;132;113m \033[48;2;182;135;115m \033[48;2;193;145;124m \033[48;2;200;152;131m \033[48;2;201;150;129m \033[48;2;203;154;133m \033[48;2;210;159;138m \033[48;2;209;158;135m \033[48;2;202;148;124m \033[48;2;200;143;121m \033[48;2;204;146;123m \033[48;2;205;148;125m \033[48;2;203;147;124m \033[48;2;205;148;126m \033[48;2;202;145;123m \033[48;2;198;141;121m \033[48;2;194;138;118m \033[48;2;183;129;109m \033[48;2;171;119;99m \033[48;2;164;113;94m \033[48;2;157;107;91m \033[48;2;145;99;86m \033[48;2;129;89;81m \033[48;2;117;80;77m \033[48;2;71;48;45m \033[48;2;45;33;35m \033[48;2;35;30;36m \033[48;2;31;29;34m \033[48;2;32;27;34m \033[48;2;57;55;60m \033[48;2;57;55;58m \033[48;2;56;54;57m \033[48;2;56;54;56m \033[48;2;53;53;53m \033[48;2;53;51;54m \033[48;2;51;50;52m \033[48;2;52;47;53m \033[48;2;50;45;51m \033[48;2;50;45;51m \033[48;2;48;43;50m \033[48;2;47;42;48m \033[48;2;46;41;47m \033[48;2;46;41;47m \033[48;2;46;41;47m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;47;42;48m \033[48;2;46;41;47m \033[48;2;45;40;46m \033[48;2;45;39;45m \033[48;2;44;39;45m \033[48;2;43;40;44m \033[48;2;43;40;44m \033[48;2;44;42;43m \033[48;2;46;43;44m \033[48;2;45;43;42m \033[48;2;46;45;43m \033[48;2;47;45;41m \033[48;2;46;45;41m \033[48;2;45;43;39m \033[m");
$display("\033[48;2;87;85;88m \033[48;2;90;88;91m \033[48;2;98;96;99m \033[48;2;95;93;96m \033[48;2;95;93;94m \033[48;2;94;91;93m \033[48;2;93;93;93m \033[48;2;92;92;92m \033[48;2;89;89;89m \033[48;2;88;88;88m \033[48;2;88;88;88m \033[48;2;91;88;92m \033[48;2;91;88;92m \033[48;2;90;88;88m \033[48;2;90;88;89m \033[48;2;91;89;90m \033[48;2;94;92;94m \033[48;2;88;86;87m \033[48;2;86;83;85m \033[48;2;86;84;85m \033[48;2;83;81;84m \033[48;2;79;77;78m \033[48;2;72;71;69m \033[48;2;68;67;63m \033[48;2;65;65;63m \033[48;2;61;61;59m \033[48;2;60;59;57m \033[48;2;55;55;53m \033[48;2;55;54;52m \033[48;2;55;55;53m \033[48;2;89;83;90m \033[48;2;62;57;63m \033[48;2;38;31;38m \033[48;2;61;49;52m \033[48;2;89;73;73m \033[48;2;97;75;72m \033[48;2;102;75;67m \033[48;2;105;75;66m \033[48;2;110;77;66m \033[48;2;112;78;65m \033[48;2;120;84;71m \033[48;2;121;82;69m \033[48;2;120;78;62m \033[48;2;110;66;51m \033[48;2;123;78;58m \033[48;2;153;106;87m \033[48;2;173;126;107m \033[48;2;189;142;124m \033[48;2;225;181;162m \033[48;2;229;186;167m \033[48;2;239;196;177m \033[48;2;245;206;185m \033[48;2;236;195;175m \033[48;2;210;168;146m \033[48;2;236;191;169m \033[48;2;251;205;182m \033[48;2;255;211;190m \033[48;2;249;204;183m \033[48;2;242;197;175m \033[48;2;220;176;155m \033[48;2;213;164;142m \033[48;2;200;153;130m \033[48;2;188;136;118m \033[48;2;181;130;111m \033[48;2;174;123;106m \033[48;2;158;109;94m \033[48;2;144;98;85m \033[48;2;136;96;86m \033[48;2;121;85;76m \033[48;2;79;57;54m \033[48;2;42;29;32m \033[48;2;33;28;34m \033[48;2;30;28;33m \033[48;2;36;32;38m \033[48;2;50;48;53m \033[48;2;50;48;51m \033[48;2;51;49;52m \033[48;2;51;49;51m \033[48;2;49;49;49m \033[48;2;49;47;50m \033[48;2;47;45;48m \033[48;2;47;42;48m \033[48;2;44;38;44m \033[48;2;45;40;46m \033[48;2;45;40;46m \033[48;2;44;39;45m \033[48;2;43;38;44m \033[48;2;44;39;45m \033[48;2;44;39;45m \033[48;2;44;39;45m \033[48;2;45;40;46m \033[48;2;46;40;47m \033[48;2;47;40;47m \033[48;2;47;40;47m \033[48;2;46;39;46m \033[48;2;45;38;45m \033[48;2;46;39;46m \033[48;2;46;39;46m \033[48;2;46;39;46m \033[48;2;46;39;46m \033[48;2;46;40;46m \033[48;2;46;40;44m \033[48;2;45;39;43m \033[48;2;45;39;41m \033[48;2;45;39;41m \033[48;2;44;38;40m \033[48;2;44;38;40m \033[48;2;45;39;39m \033[48;2;46;40;40m \033[48;2;46;42;41m \033[m");
$display("\033[48;2;86;85;87m \033[48;2;87;85;88m \033[48;2;86;84;85m \033[48;2;85;83;86m \033[48;2;83;81;84m \033[48;2;81;79;83m \033[48;2;80;78;81m \033[48;2;78;76;79m \033[48;2;76;74;77m \033[48;2;75;73;76m \033[48;2;74;72;75m \033[48;2;72;71;76m \033[48;2;71;70;75m \033[48;2;69;68;73m \033[48;2;69;68;73m \033[48;2;69;68;73m \033[48;2;66;65;70m \033[48;2;62;61;66m \033[48;2;60;59;64m \033[48;2;57;56;61m \033[48;2;55;54;60m \033[48;2;54;53;59m \033[48;2;52;49;56m \033[48;2;51;48;55m \033[48;2;49;46;53m \033[48;2;48;46;51m \033[48;2;51;46;52m \033[48;2;52;46;50m \033[48;2;53;47;51m \033[48;2;51;47;47m \033[48;2;60;54;56m \033[48;2;55;47;48m \033[48;2;41;32;34m \033[48;2;85;66;63m \033[48;2;95;75;69m \033[48;2;96;73;63m \033[48;2;90;64;51m \033[48;2;84;54;43m \033[48;2;91;57;47m \033[48;2;92;56;44m \033[48;2;91;55;43m \033[48;2;92;55;41m \033[48;2;94;55;38m \033[48;2;104;67;48m \033[48;2;103;67;45m \033[48;2;110;68;46m \033[48;2;123;77;55m \033[48;2;154;103;82m \033[48;2;182;134;112m \033[48;2;214;168;145m \033[48;2;213;167;144m \033[48;2;213;168;142m \033[48;2;210;164;140m \033[48;2;210;164;140m \033[48;2;218;172;150m \033[48;2;215;171;147m \033[48;2;212;171;146m \033[48;2;197;152;129m \033[48;2;168;122;99m \033[48;2;142;94;72m \033[48;2;134;85;63m \033[48;2;123;78;55m \033[48;2;111;70;48m \033[48;2;116;72;52m \033[48;2;108;62;43m \033[48;2;121;74;55m \033[48;2;122;76;61m \033[48;2;133;92;79m \033[48;2;132;97;85m \033[48;2;88;67;60m \033[48;2;44;32;31m \033[48;2;37;33;34m \033[48;2;36;33;36m \033[48;2;48;42;44m \033[48;2;52;47;51m \033[48;2;52;47;51m \033[48;2;49;44;48m \033[48;2;47;42;46m \033[48;2;45;40;44m \033[48;2;45;40;44m \033[48;2;45;40;44m \033[48;2;41;36;40m \033[48;2;43;38;43m \033[48;2;40;38;43m \033[48;2;40;38;43m \033[48;2;41;39;43m \033[48;2;41;39;42m \033[48;2;41;40;42m \033[48;2;40;38;41m \033[48;2;37;34;35m \033[48;2;27;23;22m \033[48;2;17;12;12m \033[48;2;19;11;9m \033[48;2;21;13;11m \033[48;2;26;18;16m \033[48;2;37;29;27m \033[48;2;37;27;26m \033[48;2;35;25;24m \033[48;2;33;23;22m \033[48;2;33;23;22m \033[48;2;32;22;21m \033[48;2;28;18;17m \033[48;2;24;15;13m \033[48;2;25;15;14m \033[48;2;25;15;14m \033[48;2;26;16;17m \033[48;2;28;18;19m \033[48;2;36;26;27m \033[48;2;37;27;28m \033[48;2;43;33;35m \033[m");
$display("\033[48;2;84;84;86m \033[48;2;84;82;85m \033[48;2;81;79;82m \033[48;2;77;75;80m \033[48;2;75;73;78m \033[48;2;70;69;75m \033[48;2;69;67;71m \033[48;2;66;64;69m \033[48;2;61;59;64m \033[48;2;60;58;63m \033[48;2;58;56;61m \033[48;2;54;53;58m \033[48;2;52;51;56m \033[48;2;53;52;57m \033[48;2;54;53;58m \033[48;2;54;54;56m \033[48;2;51;51;53m \033[48;2;47;47;49m \033[48;2;44;44;46m \033[48;2;43;43;43m \033[48;2;43;42;48m \033[48;2;48;47;53m \033[48;2;43;40;47m \033[48;2;39;36;43m \033[48;2;35;32;39m \033[48;2;32;30;35m \033[48;2;30;25;31m \033[48;2;31;25;29m \033[48;2;93;86;90m \033[48;2;91;80;84m \033[48;2;54;40;40m \033[48;2;53;35;34m \033[48;2;54;34;30m \033[48;2;96;71;65m \033[48;2;101;74;65m \033[48;2;101;71;63m \033[48;2;106;73;64m \033[48;2;109;75;66m \033[48;2;116;82;72m \033[48;2;142;105;94m \033[48;2;166;130;118m \033[48;2;187;150;137m \033[48;2;194;155;139m \033[48;2;195;158;140m \033[48;2;178;141;123m \033[48;2;146;104;85m \033[48;2;107;62;41m \033[48;2;118;70;48m \033[48;2;137;86;65m \033[48;2;167;116;95m \033[48;2;194;142;121m \033[48;2;204;155;130m \033[48;2;206;156;133m \033[48;2;213;163;140m \033[48;2;219;169;147m \033[48;2;216;165;144m \033[48;2;202;151;130m \033[48;2;170;118;97m \033[48;2;148;97;76m \033[48;2;118;67;46m \033[48;2;116;67;45m \033[48;2;117;72;49m \033[48;2;121;79;57m \033[48;2;135;92;71m \033[48;2;135;90;71m \033[48;2;135;88;70m \033[48;2;122;76;61m \033[48;2;106;64;51m \033[48;2;134;99;87m \033[48;2;100;78;74m \033[48;2;44;31;31m \033[48;2;36;30;34m \033[48;2;43;40;45m \033[48;2;56;50;54m \033[48;2;54;49;55m \033[48;2;52;47;53m \033[48;2;51;46;52m \033[48;2;47;42;48m \033[48;2;43;38;42m \033[48;2;43;38;42m \033[48;2;43;38;42m \033[48;2;42;37;41m \033[48;2;42;37;41m \033[48;2;41;36;42m \033[48;2;40;35;39m \033[48;2;42;38;39m \033[48;2;36;32;33m \033[48;2;22;18;19m \033[48;2;18;14;13m \033[48;2;14;8;9m \033[48;2;17;12;9m \033[48;2;28;22;19m \033[48;2;39;31;29m \033[48;2;38;30;28m \033[48;2;38;30;28m \033[48;2;38;30;28m \033[48;2;39;29;28m \033[48;2;39;29;28m \033[48;2;38;28;27m \033[48;2;37;27;26m \033[48;2;37;27;26m \033[48;2;37;27;26m \033[48;2;37;27;26m \033[48;2;37;27;26m \033[48;2;37;27;26m \033[48;2;38;28;27m \033[48;2;38;28;27m \033[48;2;38;28;27m \033[48;2;38;28;27m \033[48;2;56;46;46m \033[m");
$display("\033[48;2;89;86;95m \033[48;2;83;79;93m \033[48;2;73;70;79m \033[48;2;66;63;72m \033[48;2;61;58;65m \033[48;2;56;53;60m \033[48;2;52;49;56m \033[48;2;52;49;56m \033[48;2;51;48;55m \033[48;2;50;47;54m \033[48;2;47;45;52m \033[48;2;41;40;46m \033[48;2;38;37;43m \033[48;2;35;34;40m \033[48;2;34;33;39m \033[48;2;31;31;37m \033[48;2;31;30;36m \033[48;2;48;47;53m \033[48;2;53;52;59m \033[48;2;61;60;66m \033[48;2;40;39;48m \033[48;2;32;30;40m \033[48;2;39;37;46m \033[48;2;29;28;36m \033[48;2;35;28;39m \033[48;2;32;29;38m \033[48;2;40;33;40m \033[48;2;69;52;55m \033[48;2;101;72;76m \033[48;2;104;74;77m \033[48;2;73;49;50m \033[48;2;59;33;32m \033[48;2;68;40;37m \033[48;2;102;69;64m \033[48;2;107;69;61m \033[48;2;122;84;73m \033[48;2;140;103;93m \033[48;2;137;101;91m \033[48;2;127;87;77m \033[48;2;103;64;54m \033[48;2;78;40;31m \033[48;2;67;30;21m \033[48;2;60;26;17m \033[48;2;69;38;24m \033[48;2;95;60;44m \033[48;2;153;115;96m \033[48;2;143;96;77m \033[48;2;144;94;77m \033[48;2;118;65;46m \033[48;2;107;52;34m \033[48;2;174;119;97m \033[48;2;217;166;141m \033[48;2;230;182;159m \033[48;2;239;191;168m \033[48;2;207;157;135m \033[48;2;144;89;69m \033[48;2;151;93;76m \033[48;2;165;112;92m \033[48;2;177;127;110m \033[48;2;185;137;124m \033[48;2;207;164;148m \033[48;2;209;171;152m \033[48;2;214;176;155m \033[48;2;203;162;141m \033[48;2;201;158;137m \033[48;2;190;143;127m \033[48;2;167;120;103m \033[48;2;141;99;85m \033[48;2;128;93;82m \033[48;2;108;86;80m \033[48;2;45;30;29m \033[48;2;36;26;30m \033[48;2;51;43;47m \033[48;2;56;48;52m \033[48;2;54;49;56m \033[48;2;52;47;54m \033[48;2;47;42;49m \033[48;2;45;40;47m \033[48;2;42;36;40m \033[48;2;42;36;40m \033[48;2;42;36;38m \033[48;2;42;36;38m \033[48;2;43;37;39m \033[48;2;43;39;40m \033[48;2;46;42;43m \033[48;2;26;21;25m \033[48;2;17;12;17m \033[48;2;15;14;12m \033[48;2;16;11;15m \033[48;2;21;16;20m \033[48;2;35;26;28m \033[48;2;43;33;32m \033[48;2;44;32;32m \033[48;2;43;33;32m \033[48;2;41;32;30m \033[48;2;42;34;31m \033[48;2;41;34;27m \033[48;2;41;33;28m \033[48;2;39;30;29m \033[48;2;36;27;28m \033[48;2;35;26;29m \033[48;2;33;26;31m \033[48;2;34;27;31m \033[48;2;41;28;26m \033[48;2;36;26;24m \033[48;2;40;30;26m \033[48;2;43;31;33m \033[48;2;46;33;40m \033[48;2;46;35;43m \033[48;2;61;49;57m \033[m");
$display("\033[48;2;39;36;44m \033[48;2;48;43;58m \033[48;2;67;65;76m \033[48;2;43;40;51m \033[48;2;34;32;41m \033[48;2;27;24;33m \033[48;2;18;15;22m \033[48;2;8;5;12m \033[48;2;6;3;10m \033[48;2;7;4;11m \033[48;2;8;5;12m \033[48;2;8;5;12m \033[48;2;11;8;15m \033[48;2;23;20;27m \033[48;2;27;24;31m \033[48;2;19;16;23m \033[48;2;18;15;22m \033[48;2;14;11;18m \033[48;2;14;11;18m \033[48;2;12;9;15m \033[48;2;15;12;21m \033[48;2;13;10;19m \033[48;2;13;9;18m \033[48;2;17;14;24m \033[48;2;21;19;25m \033[48;2;23;19;26m \033[48;2;44;34;40m \033[48;2;89;67;69m \033[48;2;101;65;70m \033[48;2;107;67;70m \033[48;2;67;36;32m \033[48;2;58;32;23m \033[48;2;92;65;53m \033[48;2;109;75;62m \033[48;2;124;86;68m \033[48;2;137;94;77m \033[48;2;132;89;72m \033[48;2;117;73;58m \033[48;2;113;70;54m \033[48;2;150;108;94m \033[48;2;162;121;107m \033[48;2;155;115;101m \033[48;2;113;75;64m \033[48;2;99;63;51m \033[48;2;146;110;96m \033[48;2;205;167;152m \033[48;2;185;141;126m \033[48;2;179;127;111m \033[48;2;190;137;120m \033[48;2;143;88;69m \033[48;2;184;129;108m \033[48;2;210;159;134m \033[48;2;229;182;156m \033[48;2;226;178;154m \033[48;2;197;146;124m \033[48;2;193;137;118m \033[48;2;174;116;100m \033[48;2;169;114;94m \033[48;2;188;139;122m \033[48;2;102;56;41m \033[48;2;97;58;41m \033[48;2;97;61;41m \033[48;2;117;79;60m \033[48;2;141;97;78m \033[48;2;161;113;96m \033[48;2;182;132;118m \033[48;2;175;127;112m \033[48;2;147;103;90m \033[48;2;131;94;84m \033[48;2;97;70;67m \033[48;2;48;27;29m \033[48;2;38;24;31m \033[48;2;53;40;49m \033[48;2;58;47;53m \033[48;2;51;44;51m \033[48;2;48;41;48m \033[48;2;45;38;45m \033[48;2;44;37;44m \033[48;2;40;35;39m \033[48;2;40;35;39m \033[48;2;42;38;39m \033[48;2;44;40;41m \033[48;2;46;42;43m \033[48;2;39;35;37m \033[48;2;23;19;19m \033[48;2;18;13;17m \033[48;2;17;12;16m \033[48;2;14;11;11m \033[48;2;20;13;20m \033[48;2;35;26;34m \033[48;2;39;28;32m \033[48;2;65;50;51m \033[48;2;68;54;51m \033[48;2;74;55;50m \033[48;2;80;58;51m \033[48;2;94;69;60m \033[48;2;120;94;81m \033[48;2;124;98;84m \033[48;2;135;110;94m \033[48;2;157;132;117m \033[48;2;163;138;119m \033[48;2;153;130;97m \033[48;2;148;128;93m \033[48;2;124;105;96m \033[48;2;103;83;82m \033[48;2;79;63;64m \033[48;2;70;54;53m \033[48;2;61;45;45m \033[48;2;68;53;58m \033[48;2;66;53;63m \033[m");
$display("\033[48;2;53;52;61m \033[48;2;54;52;65m \033[48;2;23;19;33m \033[48;2;6;3;14m \033[48;2;7;4;15m \033[48;2;5;2;13m \033[48;2;6;1;8m \033[48;2;6;1;8m \033[48;2;7;1;8m \033[48;2;8;3;10m \033[48;2;8;3;10m \033[48;2;8;5;12m \033[48;2;11;9;16m \033[48;2;20;19;25m \033[48;2;19;18;24m \033[48;2;15;14;20m \033[48;2;14;11;18m \033[48;2;14;11;18m \033[48;2;13;10;17m \033[48;2;11;8;15m \033[48;2;11;8;15m \033[48;2;11;8;15m \033[48;2;11;8;15m \033[48;2;12;9;16m \033[48;2;13;12;17m \033[48;2;16;14;19m \033[48;2;20;12;14m \033[48;2;88;65;67m \033[48;2;99;63;63m \033[48;2;117;78;77m \033[48;2;87;53;45m \033[48;2;69;33;21m \033[48;2;109;71;55m \033[48;2;123;82;63m \033[48;2;140;98;74m \033[48;2;156;108;85m \033[48;2;161;111;90m \033[48;2;163;112;93m \033[48;2;167;115;94m \033[48;2;169;117;96m \033[48;2;170;115;95m \033[48;2;180;123;104m \033[48;2;180;125;104m \033[48;2;170;118;96m \033[48;2;174;122;101m \033[48;2;195;143;122m \033[48;2;225;173;152m \033[48;2;201;152;131m \033[48;2;153;101;80m \033[48;2;172;117;96m \033[48;2;201;147;126m \033[48;2;227;175;153m \033[48;2;234;187;164m \033[48;2;228;183;159m \033[48;2;206;156;135m \033[48;2;213;160;142m \033[48;2;184;133;112m \033[48;2;190;142;122m \033[48;2;205;161;142m \033[48;2;159;119;100m \033[48;2;142;100;84m \033[48;2;157;118;100m \033[48;2;196;156;138m \033[48;2;176;132;111m \033[48;2;155;103;87m \033[48;2;171;116;101m \033[48;2;171;119;105m \033[48;2;162;114;104m \033[48;2;136;94;87m \033[48;2;95;65;61m \033[48;2;55;25;23m \033[48;2;54;23;26m \033[48;2;91;62;66m \033[48;2;101;76;79m \033[48;2;67;45;52m \033[48;2;51;38;45m \033[48;2;45;39;43m \033[48;2;47;38;41m \033[48;2;46;39;45m \033[48;2;47;41;45m \033[48;2;49;44;48m \033[48;2;52;48;49m \033[48;2;48;44;45m \033[48;2;20;16;17m \033[48;2;20;17;17m \033[48;2;16;11;15m \033[48;2;16;11;16m \033[48;2;17;12;18m \033[48;2;24;19;25m \033[48;2;32;24;32m \033[48;2;51;38;46m \033[48;2;68;51;56m \033[48;2;94;71;68m \033[48;2;103;78;88m \033[48;2;69;55;86m \033[48;2;64;57;90m \033[48;2;70;58;93m \033[48;2;70;58;93m \033[48;2;74;63;97m \033[48;2;73;62;96m \033[48;2;82;68;98m \033[48;2;121;97;103m \033[48;2;79;67;75m \033[48;2;62;65;104m \033[48;2;61;63;109m \033[48;2;57;59;102m \033[48;2;58;57;96m \033[48;2;63;53;87m \033[48;2;67;54;76m \033[48;2;69;54;69m \033[m");
$display("\033[48;2;51;52;60m \033[48;2;51;51;63m \033[48;2;11;8;19m \033[48;2;4;1;12m \033[48;2;4;1;10m \033[48;2;3;0;9m \033[48;2;3;1;6m \033[48;2;3;1;6m \033[48;2;4;2;7m \033[48;2;6;4;9m \033[48;2;6;4;9m \033[48;2;8;7;13m \033[48;2;17;16;22m \033[48;2;19;20;25m \033[48;2;17;19;24m \033[48;2;13;15;20m \033[48;2;12;13;17m \033[48;2;11;10;16m \033[48;2;9;8;14m \033[48;2;8;7;13m \033[48;2;8;6;11m \033[48;2;8;6;11m \033[48;2;10;8;13m \033[48;2;11;9;14m \033[48;2;14;12;17m \033[48;2;16;14;19m \033[48;2;20;12;16m \033[48;2;56;33;35m \033[48;2;98;62;62m \033[48;2;107;68;63m \033[48;2;101;61;54m \033[48;2;103;61;48m \033[48;2;121;77;62m \033[48;2;127;80;62m \033[48;2;138;90;68m \033[48;2;163;113;86m \033[48;2;178;125;98m \033[48;2;189;133;108m \033[48;2;192;136;110m \033[48;2;198;142;117m \033[48;2;203;147;121m \033[48;2;203;148;120m \033[48;2;203;149;121m \033[48;2;207;153;124m \033[48;2;211;156;130m \033[48;2;211;157;131m \033[48;2;191;137;111m \033[48;2;162;106;83m \033[48;2;168;107;86m \033[48;2;191;130;108m \033[48;2;218;160;140m \033[48;2;235;183;161m \033[48;2;238;189;167m \033[48;2;235;188;165m \033[48;2;215;165;144m \033[48;2;212;159;138m \033[48;2;219;168;147m \033[48;2;219;171;149m \033[48;2;200;153;133m \033[48;2;180;133;113m \033[48;2;183;131;115m \033[48;2;192;141;121m \033[48;2;207;156;135m \033[48;2;206;153;131m \033[48;2;206;154;128m \033[48;2;191;137;111m \033[48;2;189;135;111m \033[48;2;182;129;111m \033[48;2;146;98;85m \033[48;2;91;49;39m \033[48;2;82;35;29m \033[48;2;122;73;69m \033[48;2;118;71;68m \033[48;2;116;75;74m \033[48;2;93;63;65m \033[48;2;50;35;38m \033[48;2;48;39;42m \033[48;2;48;39;41m \033[48;2;46;40;44m \033[48;2;46;40;44m \033[48;2;49;45;46m \033[48;2;57;53;53m \033[48;2;27;23;21m \033[48;2;21;17;18m \033[48;2;18;14;15m \033[48;2;16;11;15m \033[48;2;16;11;15m \033[48;2;15;10;16m \033[48;2;27;22;28m \033[48;2;31;24;31m \033[48;2;49;38;46m \033[48;2;66;50;55m \033[48;2;117;95;88m \033[48;2;86;59;67m \033[48;2;69;56;95m \033[48;2;64;59;100m \033[48;2;60;59;98m \033[48;2;61;60;98m \033[48;2;63;62;98m \033[48;2;71;70;103m \033[48;2;83;80;109m \033[48;2;158;137;138m \033[48;2;69;55;62m \033[48;2;64;67;104m \033[48;2;63;67;106m \033[48;2;56;60;101m \033[48;2;56;57;98m \033[48;2;62;54;91m \033[48;2;69;55;79m \033[48;2;72;56;68m \033[m");
$display("\033[48;2;51;54;61m \033[48;2;50;50;62m \033[48;2;4;1;10m \033[48;2;5;2;11m \033[48;2;4;1;8m \033[48;2;3;0;7m \033[48;2;2;1;7m \033[48;2;2;1;7m \033[48;2;2;1;7m \033[48;2;5;4;10m \033[48;2;6;5;11m \033[48;2;15;15;20m \033[48;2;18;19;24m \033[48;2;14;17;22m \033[48;2;13;16;21m \033[48;2;8;12;15m \033[48;2;5;9;12m \033[48;2;7;8;12m \033[48;2;6;7;12m \033[48;2;6;5;10m \033[48;2;7;4;11m \033[48;2;7;4;11m \033[48;2;8;5;12m \033[48;2;9;6;13m \033[48;2;10;8;13m \033[48;2;11;9;14m \033[48;2;19;11;14m \033[48;2;55;32;34m \033[48;2;96;62;62m \033[48;2;96;55;49m \033[48;2;128;79;72m \033[48;2;123;72;59m \033[48;2;129;78;63m \033[48;2;131;79;62m \033[48;2;138;87;65m \033[48;2;166;111;81m \033[48;2;183;125;95m \033[48;2;193;134;104m \033[48;2;203;144;110m \033[48;2;211;155;120m \033[48;2;213;157;122m \033[48;2;213;161;124m \033[48;2;214;160;124m \033[48;2;216;162;128m \033[48;2;218;165;130m \033[48;2;209;155;124m \033[48;2;180;125;94m \033[48;2;164;109;78m \033[48;2;172;116;89m \033[48;2;207;151;125m \033[48;2;222;172;148m \033[48;2;238;185;163m \033[48;2;244;196;173m \033[48;2;245;199;176m \033[48;2;230;180;159m \033[48;2;218;167;146m \033[48;2;222;176;152m \033[48;2;235;189;165m \033[48;2;238;190;168m \033[48;2;232;184;162m \033[48;2;227;181;157m \033[48;2;233;183;157m \033[48;2;224;170;144m \033[48;2;225;174;145m \033[48;2;217;169;138m \033[48;2;214;160;131m \033[48;2;202;144;120m \033[48;2;192;135;117m \033[48;2;154;96;86m \033[48;2;96;49;40m \033[48;2;125;75;67m \033[48;2;152;98;96m \033[48;2;121;71;69m \033[48;2;133;88;84m \033[48;2;100;63;61m \033[48;2;60;38;40m \033[48;2;51;41;42m \033[48;2;50;41;42m \033[48;2;50;44;46m \033[48;2;50;44;46m \033[48;2;57;53;52m \033[48;2;56;52;50m \033[48;2;24;20;19m \033[48;2;19;15;16m \033[48;2;19;15;16m \033[48;2;16;11;15m \033[48;2;14;9;13m \033[48;2;16;11;17m \033[48;2;28;23;29m \033[48;2;32;25;32m \033[48;2;49;37;45m \033[48;2;65;48;52m \033[48;2;163;140;131m \033[48;2;61;35;45m \033[48;2;57;43;84m \033[48;2;52;46;90m \033[48;2;48;47;91m \033[48;2;49;48;90m \033[48;2;50;49;90m \033[48;2;51;51;89m \033[48;2;53;52;84m \033[48;2;175;156;160m \033[48;2;56;45;55m \033[48;2;51;56;95m \033[48;2;51;55;98m \033[48;2;47;55;92m \033[48;2;51;52;98m \033[48;2;57;50;92m \033[48;2;66;55;80m \033[48;2;73;59;67m \033[m");
$display("\033[48;2;53;54;59m \033[48;2;49;49;57m \033[48;2;2;1;9m \033[48;2;2;1;9m \033[48;2;1;0;8m \033[48;2;1;0;8m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;4;3;8m \033[48;2;13;12;17m \033[48;2;21;21;27m \033[48;2;17;18;23m \033[48;2;16;18;23m \033[48;2;12;15;20m \033[48;2;9;10;15m \033[48;2;9;8;14m \033[48;2;7;6;12m \033[48;2;7;6;12m \033[48;2;7;5;10m \033[48;2;6;4;9m \033[48;2;6;4;9m \033[48;2;7;5;10m \033[48;2;9;7;11m \033[48;2;9;7;10m \033[48;2;11;9;14m \033[48;2;17;6;11m \033[48;2;80;54;57m \033[48;2;100;65;62m \033[48;2;115;74;68m \033[48;2;109;60;52m \033[48;2;124;72;59m \033[48;2;130;79;64m \033[48;2;144;93;76m \033[48;2;145;89;70m \033[48;2;164;106;81m \033[48;2;184;123;93m \033[48;2;195;135;101m \033[48;2;207;150;115m \033[48;2;213;159;123m \033[48;2;219;165;128m \033[48;2;222;170;133m \033[48;2;224;173;133m \033[48;2;227;175;138m \033[48;2;227;173;139m \033[48;2;216;160;130m \033[48;2;173;118;86m \033[48;2;168;113;83m \033[48;2;198;143;116m \033[48;2;211;159;134m \033[48;2;232;182;157m \033[48;2;253;211;187m \033[48;2;255;222;198m \033[48;2;245;217;193m \033[48;2;241;204;183m \033[48;2;234;188;170m \033[48;2;230;185;162m \033[48;2;242;196;174m \033[48;2;248;203;180m \033[48;2;247;203;181m \033[48;2;245;196;174m \033[48;2;236;190;163m \033[48;2;234;184;153m \033[48;2;233;182;150m \033[48;2;233;180;149m \033[48;2;219;168;139m \033[48;2;205;151;126m \033[48;2;194;138;119m \033[48;2;161;104;85m \033[48;2;123;71;58m \033[48;2;165;111;100m \033[48;2;167;112;106m \033[48;2;141;90;88m \033[48;2;133;90;88m \033[48;2;70;40;40m \033[48;2;62;43;45m \033[48;2;54;45;48m \033[48;2;55;46;49m \033[48;2;54;48;50m \033[48;2;54;48;50m \033[48;2;58;52;52m \033[48;2;60;54;54m \033[48;2;24;18;18m \033[48;2;19;14;18m \033[48;2;19;14;19m \033[48;2;16;11;17m \033[48;2;13;8;14m \033[48;2;16;11;18m \033[48;2;31;26;33m \033[48;2;33;27;35m \033[48;2;44;30;40m \033[48;2;70;50;58m \033[48;2;182;159;145m \033[48;2;77;53;60m \033[48;2;54;46;81m \033[48;2;46;43;88m \033[48;2;44;45;92m \033[48;2;42;43;93m \033[48;2;41;43;92m \033[48;2;41;43;91m \033[48;2;42;44;83m \033[48;2;178;162;157m \033[48;2;51;40;65m \033[48;2;38;45;88m \033[48;2;41;45;92m \033[48;2;40;45;92m \033[48;2;42;44;92m \033[48;2;48;43;84m \033[48;2;65;54;78m \033[48;2;75;59;69m \033[m");
$display("\033[48;2;54;55;59m \033[48;2;39;39;46m \033[48;2;1;0;8m \033[48;2;3;2;10m \033[48;2;2;1;9m \033[48;2;1;0;8m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;2;1;6m \033[48;2;8;7;11m \033[48;2;21;20;24m \033[48;2;18;19;24m \033[48;2;19;20;25m \033[48;2;15;17;22m \033[48;2;8;10;16m \033[48;2;10;10;16m \033[48;2;7;5;12m \033[48;2;5;4;10m \033[48;2;5;3;10m \033[48;2;6;4;9m \033[48;2;6;4;7m \033[48;2;6;4;7m \033[48;2;6;4;7m \033[48;2;8;6;9m \033[48;2;8;6;7m \033[48;2;9;7;10m \033[48;2;13;4;4m \033[48;2;106;80;79m \033[48;2;119;84;80m \033[48;2;121;80;74m \033[48;2;123;74;66m \033[48;2;108;57;44m \033[48;2;124;72;57m \033[48;2;154;103;85m \033[48;2;159;103;85m \033[48;2;164;107;83m \033[48;2;177;116;85m \033[48;2;195;134;100m \033[48;2;205;146;112m \033[48;2;217;158;124m \033[48;2;219;163;128m \033[48;2;226;171;135m \033[48;2;230;176;139m \033[48;2;235;181;145m \033[48;2;243;187;154m \033[48;2;193;137;107m \033[48;2;187;127;98m \033[48;2;185;124;99m \033[48;2;182;121;100m \033[48;2;185;128;107m \033[48;2;209;153;133m \033[48;2;239;193;170m \033[48;2;241;199;177m \033[48;2;237;197;177m \033[48;2;241;198;180m \033[48;2;246;197;181m \033[48;2;236;188;170m \033[48;2;234;184;168m \033[48;2;231;184;166m \033[48;2;244;197;179m \033[48;2;254;209;185m \033[48;2;255;209;182m \033[48;2;242;196;163m \033[48;2;237;186;155m \033[48;2;231;180;149m \033[48;2;224;175;142m \033[48;2;206;155;126m \033[48;2;191;137;114m \033[48;2;158;103;82m \033[48;2;180;122;109m \033[48;2;183;125;114m \033[48;2;171;117;109m \033[48;2;139;90;86m \033[48;2;87;48;44m \033[48;2;63;40;43m \033[48;2;55;44;48m \033[48;2;53;47;49m \033[48;2;56;47;48m \033[48;2;55;49;49m \033[48;2;58;52;54m \033[48;2;57;51;55m \033[48;2;56;49;56m \033[48;2;20;13;20m \033[48;2;19;14;20m \033[48;2;18;13;19m \033[48;2;14;9;16m \033[48;2;10;6;13m \033[48;2;13;8;16m \033[48;2;30;25;32m \033[48;2;36;29;37m \033[48;2;38;26;36m \033[48;2;78;57;65m \033[48;2;161;133;117m \033[48;2;82;58;65m \033[48;2;48;42;79m \033[48;2;41;42;90m \033[48;2;41;41;91m \033[48;2;37;40;90m \033[48;2;32;39;88m \033[48;2;29;40;86m \033[48;2;35;43;81m \033[48;2;144;131;125m \033[48;2;42;36;63m \033[48;2;27;39;81m \033[48;2;29;37;83m \033[48;2;26;35;82m \033[48;2;28;34;88m \033[48;2;36;37;83m \033[48;2;67;54;80m \033[48;2;74;53;62m \033[m");
$display("\033[48;2;52;53;58m \033[48;2;30;29;37m \033[48;2;0;0;7m \033[48;2;3;2;8m \033[48;2;2;1;7m \033[48;2;1;0;5m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;3;2;9m \033[48;2;20;19;26m \033[48;2;22;22;27m \033[48;2;17;20;25m \033[48;2;18;21;26m \033[48;2;17;19;24m \033[48;2;10;13;18m \033[48;2;6;11;15m \033[48;2;2;5;10m \033[48;2;4;5;10m \033[48;2;5;4;10m \033[48;2;5;4;9m \033[48;2;6;4;7m \033[48;2;6;4;7m \033[48;2;6;4;7m \033[48;2;8;6;9m \033[48;2;9;7;10m \033[48;2;11;10;13m \033[48;2;19;10;12m \033[48;2;53;31;29m \033[48;2;112;78;74m \033[48;2;116;73;67m \033[48;2;108;61;54m \033[48;2;83;33;22m \033[48;2;118;69;51m \033[48;2;146;96;80m \033[48;2;153;98;78m \033[48;2;161;99;74m \033[48;2;170;104;74m \033[48;2;185;119;85m \033[48;2;196;132;99m \033[48;2;206;143;110m \033[48;2;218;156;120m \033[48;2;226;166;130m \033[48;2;227;170;133m \033[48;2;227;169;135m \033[48;2;198;137;105m \033[48;2;127;63;35m \033[48;2;112;46;19m \033[48;2;100;31;9m \033[48;2;94;26;6m \033[48;2;91;26;6m \033[48;2;122;58;39m \033[48;2;162;96;79m \033[48;2;152;87;70m \033[48;2;169;105;90m \033[48;2;124;64;51m \033[48;2;104;44;31m \033[48;2;139;76;61m \033[48;2;204;140;125m \033[48;2;239;175;158m \033[48;2;216;153;135m \033[48;2;227;172;151m \033[48;2;246;195;170m \033[48;2;244;194;165m \033[48;2;245;193;162m \033[48;2;243;188;157m \033[48;2;232;179;148m \033[48;2;209;156;125m \033[48;2;186;132;107m \033[48;2;174;118;99m \033[48;2;170;114;99m \033[48;2;175;115;105m \033[48;2;162;104;100m \033[48;2;144;96;93m \033[48;2;78;44;43m \033[48;2;63;43;44m \033[48;2;55;45;44m \033[48;2;53;47;49m \033[48;2;57;48;51m \033[48;2;58;52;52m \033[48;2;60;54;54m \033[48;2;60;56;57m \033[48;2;62;58;61m \033[48;2;33;28;32m \033[48;2;18;13;17m \033[48;2;19;14;21m \033[48;2;13;8;14m \033[48;2;9;4;8m \033[48;2;10;6;9m \033[48;2;21;16;22m \033[48;2;37;28;36m \033[48;2;39;24;32m \033[48;2;66;45;46m \033[48;2;118;89;82m \033[48;2;79;58;70m \033[48;2;45;37;82m \033[48;2;42;38;90m \033[48;2;41;41;86m \033[48;2;38;39;83m \033[48;2;35;38;81m \033[48;2;36;42;83m \033[48;2;63;62;94m \033[48;2;87;69;75m \033[48;2;44;23;51m \033[48;2;28;28;63m \033[48;2;28;29;62m \033[48;2;33;26;65m \033[48;2;26;23;57m \033[48;2;34;25;57m \033[48;2;67;53;72m \033[48;2;69;52;55m \033[m");
$display("\033[48;2;55;56;61m \033[48;2;17;17;25m \033[48;2;1;0;8m \033[48;2;1;0;7m \033[48;2;2;1;7m \033[48;2;1;0;5m \033[48;2;2;1;7m \033[48;2;0;0;5m \033[48;2;17;16;22m \033[48;2;29;28;34m \033[48;2;22;23;28m \033[48;2;17;21;26m \033[48;2;19;22;27m \033[48;2;12;14;20m \033[48;2;11;14;19m \033[48;2;5;8;13m \033[48;2;5;6;11m \033[48;2;4;3;9m \033[48;2;4;1;8m \033[48;2;5;0;6m \033[48;2;8;3;7m \033[48;2;9;4;8m \033[48;2;11;6;10m \033[48;2;14;9;13m \033[48;2;18;10;18m \033[48;2;19;13;15m \033[48;2;24;17;15m \033[48;2;26;16;15m \033[48;2;27;16;17m \033[48;2;23;15;12m \033[48;2;26;15;11m \033[48;2;33;15;8m \033[48;2;90;67;56m \033[48;2;135;93;74m \033[48;2;154;100;79m \033[48;2;170;104;80m \033[48;2;173;104;75m \033[48;2;174;104;72m \033[48;2;183;112;80m \033[48;2;195;127;93m \033[48;2;203;135;99m \033[48;2;212;146;111m \033[48;2;223;158;123m \033[48;2;221;156;125m \033[48;2;220;155;125m \033[48;2;218;153;125m \033[48;2;220;153;128m \033[48;2;215;147;126m \033[48;2;199;131;112m \033[48;2;187;119;102m \033[48;2;199;132;116m \033[48;2;205;143;128m \033[48;2;194;130;115m \033[48;2;229;166;151m \033[48;2;250;187;172m \033[48;2;244;181;167m \033[48;2;241;182;164m \033[48;2;242;184;163m \033[48;2;243;185;165m \033[48;2;244;187;165m \033[48;2;205;144;119m \033[48;2;230;172;145m \033[48;2;234;181;151m \033[48;2;231;178;147m \033[48;2;233;178;148m \033[48;2;224;169;139m \033[48;2;194;139;109m \033[48;2;172;116;92m \033[48;2;173;116;97m \033[48;2;186;129;118m \033[48;2;187;128;122m \033[48;2;165;112;111m \033[48;2;100;60;59m \033[48;2;72;46;46m \033[48;2;61;47;46m \033[48;2;56;46;45m \033[48;2;57;48;51m \033[48;2;59;50;53m \033[48;2;61;52;55m \033[48;2;64;55;56m \033[48;2;65;59;59m \033[48;2;64;59;56m \033[48;2;60;55;52m \033[48;2;16;12;13m \033[48;2;17;12;18m \033[48;2;15;9;14m \033[48;2;10;6;6m \033[48;2;9;4;8m \033[48;2;10;5;11m \033[48;2;31;21;30m \033[48;2;39;24;33m \033[48;2;44;22;29m \033[48;2;115;92;90m \033[48;2;112;90;88m \033[48;2;104;77;78m \033[48;2;97;75;69m \033[48;2;96;68;68m \033[48;2;89;56;63m \033[48;2;84;48;56m \033[48;2;82;43;45m \033[48;2;116;81;74m \033[48;2;200;168;137m \033[48;2;208;166;141m \033[48;2;205;160;132m \033[48;2;196;151;114m \033[48;2;193;155;114m \033[48;2;180;148;110m \033[48;2;154;131;95m \033[48;2;84;59;38m \033[48;2;64;39;34m \033[m");
$display("\033[48;2;54;55;59m \033[48;2;4;5;10m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;0;0;5m \033[48;2;0;0;4m \033[48;2;8;7;14m \033[48;2;28;27;33m \033[48;2;23;22;30m \033[48;2;22;22;30m \033[48;2;20;22;28m \033[48;2;16;19;24m \033[48;2;11;14;19m \033[48;2;8;11;16m \033[48;2;6;5;11m \033[48;2;4;3;9m \033[48;2;3;2;8m \033[48;2;4;3;9m \033[48;2;6;5;10m \033[48;2;10;5;9m \033[48;2;11;6;10m \033[48;2;12;7;11m \033[48;2;13;8;12m \033[48;2;17;11;15m \033[48;2;18;12;16m \033[48;2;21;12;17m \033[48;2;21;12;17m \033[48;2;23;12;18m \033[48;2;22;13;16m \033[48;2;24;14;13m \033[48;2;29;14;7m \033[48;2;77;54;43m \033[48;2;135;93;73m \033[48;2;161;110;89m \033[48;2;191;132;106m \033[48;2;200;137;107m \033[48;2;185;120;85m \033[48;2;186;117;84m \033[48;2;200;131;98m \033[48;2;207;138;105m \033[48;2;203;134;101m \033[48;2;207;143;108m \033[48;2;213;147;115m \033[48;2;210;143;114m \033[48;2;214;144;118m \033[48;2;217;147;122m \033[48;2;219;152;130m \033[48;2;224;159;138m \033[48;2;233;171;152m \033[48;2;244;185;167m \033[48;2;238;188;172m \033[48;2;235;182;166m \033[48;2;241;186;171m \033[48;2;245;188;173m \033[48;2;236;180;163m \033[48;2;223;166;147m \033[48;2;220;162;142m \033[48;2;233;173;154m \033[48;2;243;182;161m \033[48;2;248;182;160m \033[48;2;213;151;126m \033[48;2;232;172;146m \033[48;2;216;159;130m \033[48;2;183;127;97m \033[48;2;200;143;113m \033[48;2;200;147;116m \033[48;2;178;125;101m \033[48;2;182;128;111m \033[48;2;178;125;116m \033[48;2;177;126;122m \033[48;2;130;89;89m \033[48;2;81;54;54m \033[48;2;69;53;53m \033[48;2;65;57;55m \033[48;2;59;50;48m \033[48;2;57;48;47m \033[48;2;59;50;51m \033[48;2;62;54;51m \033[48;2;64;56;54m \033[48;2;67;59;57m \033[48;2;68;59;60m \033[48;2;68;60;61m \033[48;2;28;22;26m \033[48;2;20;14;18m \033[48;2;21;15;19m \033[48;2;12;6;10m \033[48;2;10;5;9m \033[48;2;11;5;9m \033[48;2;25;16;22m \033[48;2;36;25;31m \033[48;2;35;24;26m \033[48;2;55;46;51m \033[48;2;44;37;66m \033[48;2;34;33;80m \033[48;2;28;31;72m \033[48;2;32;32;70m \033[48;2;28;32;55m \033[48;2;28;27;52m \033[48;2;34;22;36m \033[48;2;139;117;102m \033[48;2;192;163;133m \033[48;2;146;112;84m \033[48;2;150;116;89m \033[48;2;152;120;92m \033[48;2;157;124;97m \033[48;2;162;127;100m \033[48;2;138;105;80m \033[48;2;87;60;41m \033[48;2;51;29;22m \033[m");
$display("\033[48;2;43;44;49m \033[48;2;0;0;5m \033[48;2;1;0;5m \033[48;2;1;0;5m \033[48;2;1;0;5m \033[48;2;1;0;5m \033[48;2;2;3;7m \033[48;2;23;24;29m \033[48;2;25;26;31m \033[48;2;24;24;32m \033[48;2;23;23;31m \033[48;2;24;27;32m \033[48;2;10;13;18m \033[48;2;11;14;19m \033[48;2;6;9;14m \033[48;2;5;4;9m \033[48;2;3;2;7m \033[48;2;4;3;8m \033[48;2;5;4;9m \033[48;2;7;6;11m \033[48;2;10;5;9m \033[48;2;11;6;10m \033[48;2;12;7;11m \033[48;2;13;8;12m \033[48;2;14;9;13m \033[48;2;18;13;17m \033[48;2;18;12;16m \033[48;2;19;12;16m \033[48;2;20;11;16m \033[48;2;20;11;14m \033[48;2;21;11;9m \033[48;2;26;11;3m \033[48;2;81;58;46m \033[48;2;133;95;75m \033[48;2;161;114;92m \033[48;2;196;140;113m \033[48;2;202;142;110m \033[48;2;181;121;85m \033[48;2;186;122;87m \033[48;2;196;132;97m \033[48;2;204;140;105m \033[48;2;197;133;98m \033[48;2;191;125;91m \033[48;2;191;121;91m \033[48;2;196;127;98m \033[48;2;205;133;108m \033[48;2;214;141;117m \033[48;2;221;150;130m \033[48;2;221;154;135m \033[48;2;233;169;151m \033[48;2;246;185;167m \033[48;2;244;191;173m \033[48;2;243;191;173m \033[48;2;250;197;179m \033[48;2;244;193;174m \033[48;2;235;181;163m \033[48;2;232;173;156m \033[48;2;228;167;148m \033[48;2;225;164;144m \033[48;2;231;169;148m \033[48;2;243;181;158m \033[48;2;240;180;154m \033[48;2;236;179;152m \033[48;2;222;167;137m \033[48;2;211;158;127m \033[48;2;228;175;144m \033[48;2;207;155;131m \033[48;2;135;89;74m \033[48;2;105;66;59m \033[48;2;133;96;95m \033[48;2;106;76;74m \033[48;2;79;59;58m \033[48;2;72;61;59m \033[48;2;70;61;62m \033[48;2;70;61;62m \033[48;2;65;57;55m \033[48;2;56;48;45m \033[48;2;59;51;48m \033[48;2;62;54;51m \033[48;2;64;56;54m \033[48;2;68;60;58m \033[48;2;69;60;61m \033[48;2;70;62;63m \033[48;2;50;45;49m \033[48;2;11;6;10m \033[48;2;17;12;16m \033[48;2;12;7;11m \033[48;2;9;4;8m \033[48;2;11;4;8m \033[48;2;22;13;18m \033[48;2;35;24;30m \033[48;2;39;25;31m \033[48;2;50;26;22m \033[48;2;155;114;92m \033[48;2;164;108;74m \033[48;2;169;102;71m \033[48;2;162;98;71m \033[48;2;162;100;66m \033[48;2;159;95;66m \033[48;2;160;92;61m \033[48;2;154;86;50m \033[48;2;147;79;40m \033[48;2;143;69;32m \033[48;2;142;68;28m \033[48;2;137;67;25m \033[48;2;132;64;25m \033[48;2;124;61;26m \033[48;2;109;52;24m \033[48;2;101;52;30m \033[48;2;83;38;18m \033[m");
$display("\033[48;2;19;18;23m \033[48;2;0;0;5m \033[48;2;1;1;3m \033[48;2;1;0;5m \033[48;2;1;2;6m \033[48;2;1;1;7m \033[48;2;19;21;26m \033[48;2;23;26;31m \033[48;2;21;24;31m \033[48;2;21;24;31m \033[48;2;22;25;32m \033[48;2;14;17;24m \033[48;2;13;16;21m \033[48;2;10;13;18m \033[48;2;3;7;10m \033[48;2;6;6;8m \033[48;2;6;6;8m \033[48;2;7;5;8m \033[48;2;7;5;8m \033[48;2;9;4;8m \033[48;2;9;5;9m \033[48;2;11;6;10m \033[48;2;12;7;11m \033[48;2;14;9;13m \033[48;2;14;9;13m \033[48;2;16;11;15m \033[48;2;16;11;15m \033[48;2;16;11;15m \033[48;2;16;11;15m \033[48;2;16;11;15m \033[48;2;17;11;11m \033[48;2;22;9;2m \033[48;2;87;62;52m \033[48;2;137;97;77m \033[48;2;164;119;95m \033[48;2;184;131;100m \033[48;2;187;130;97m \033[48;2;181;121;87m \033[48;2;183;119;84m \033[48;2;214;151;116m \033[48;2;213;150;115m \033[48;2;188;125;90m \033[48;2;160;96;62m \033[48;2;110;44;12m \033[48;2;122;53;24m \033[48;2;127;55;30m \033[48;2;152;80;56m \033[48;2;160;91;70m \033[48;2;169;101;82m \033[48;2;176;104;90m \033[48;2;177;105;93m \033[48;2;180;104;93m \033[48;2;187;111;101m \033[48;2;190;117;103m \033[48;2;187;113;100m \033[48;2;188;114;101m \033[48;2;163;93;79m \033[48;2;187;114;101m \033[48;2;207;136;121m \033[48;2;196;124;109m \033[48;2;213;151;128m \033[48;2;235;178;151m \033[48;2;240;183;156m \033[48;2;214;161;131m \033[48;2;244;193;162m \033[48;2;240;186;160m \033[48;2;206;156;135m \033[48;2;98;60;51m \033[48;2;82;61;59m \033[48;2;78;64;63m \033[48;2;76;64;64m \033[48;2;72;62;61m \033[48;2;71;62;63m \033[48;2;71;62;64m \033[48;2;66;63;64m \033[48;2;65;59;59m \033[48;2;55;47;44m \033[48;2;56;48;44m \033[48;2;60;52;49m \033[48;2;62;54;51m \033[48;2;67;60;57m \033[48;2;69;61;59m \033[48;2;69;61;62m \033[48;2;71;65;70m \033[48;2;22;17;21m \033[48;2;18;12;16m \033[48;2;19;13;17m \033[48;2;10;4;6m \033[48;2;7;3;4m \033[48;2;11;7;8m \033[48;2;25;15;19m \033[48;2;42;27;32m \033[48;2;48;23;28m \033[48;2;110;60;46m \033[48;2;156;83;52m \033[48;2;160;79;51m \033[48;2;159;78;49m \033[48;2;159;76;48m \033[48;2;156;76;46m \033[48;2;155;76;45m \033[48;2;156;76;46m \033[48;2;153;74;43m \033[48;2;154;73;43m \033[48;2;154;72;42m \033[48;2;157;78;47m \033[48;2;156;76;46m \033[48;2;155;80;49m \033[48;2;150;76;47m \033[48;2;144;74;46m \033[48;2;140;68;39m \033[m");
$display("\033[48;2;11;10;15m \033[48;2;1;0;5m \033[48;2;1;1;1m \033[48;2;1;1;3m \033[48;2;0;1;4m \033[48;2;10;12;15m \033[48;2;23;26;31m \033[48;2;30;33;38m \033[48;2;19;22;29m \033[48;2;20;23;30m \033[48;2;19;23;32m \033[48;2;14;14;22m \033[48;2;16;17;23m \033[48;2;9;10;15m \033[48;2;7;8;12m \033[48;2;5;5;7m \033[48;2;5;5;7m \033[48;2;6;5;7m \033[48;2;7;5;8m \033[48;2;7;5;8m \033[48;2;9;4;11m \033[48;2;11;6;12m \033[48;2;11;6;12m \033[48;2;12;7;13m \033[48;2;14;9;15m \033[48;2;15;10;17m \033[48;2;16;11;17m \033[48;2;16;11;17m \033[48;2;16;11;17m \033[48;2;13;12;17m \033[48;2;16;12;13m \033[48;2;22;11;5m \033[48;2;88;63;54m \033[48;2;135;95;77m \033[48;2;163;118;93m \033[48;2;175;125;96m \033[48;2;179;125;91m \033[48;2;174;115;82m \033[48;2;177;114;81m \033[48;2;222;162;128m \033[48;2;235;176;142m \033[48;2;237;178;144m \033[48;2;214;152;117m \033[48;2;210;147;114m \033[48;2;219;152;125m \033[48;2;229;160;134m \033[48;2;241;169;147m \033[48;2;241;174;157m \033[48;2;250;185;170m \033[48;2;248;187;174m \033[48;2;251;193;182m \033[48;2;252;196;188m \033[48;2;250;193;184m \033[48;2;250;194;184m \033[48;2;243;187;176m \033[48;2;230;170;158m \033[48;2;229;163;148m \033[48;2;224;158;141m \033[48;2;230;164;146m \033[48;2;240;175;155m \033[48;2;236;178;154m \033[48;2;249;192;165m \033[48;2;224;168;142m \033[48;2;216;162;132m \033[48;2;246;192;164m \033[48;2;220;169;146m \033[48;2;140;98;79m \033[48;2;84;56;47m \033[48;2;70;59;59m \033[48;2;74;65;68m \033[48;2;74;65;68m \033[48;2;72;66;70m \033[48;2;72;66;70m \033[48;2;71;66;69m \033[48;2;68;64;65m \033[48;2;67;62;59m \033[48;2;56;48;46m \033[48;2;57;50;46m \033[48;2;60;52;49m \033[48;2;62;54;51m \033[48;2;67;59;57m \033[48;2;67;59;57m \033[48;2;69;60;61m \033[48;2;67;61;65m \033[48;2;41;35;39m \033[48;2;15;10;14m \033[48;2;15;11;15m \033[48;2;10;5;9m \033[48;2;6;4;8m \033[48;2;8;3;7m \033[48;2;19;12;16m \033[48;2;38;25;29m \033[48;2;42;21;24m \033[48;2;66;25;17m \033[48;2;191;134;104m \033[48;2;221;154;119m \033[48;2;208;142;107m \033[48;2;172;104;69m \033[48;2;155;82;49m \033[48;2;196;122;89m \033[48;2;222;147;115m \033[48;2;191;121;87m \033[48;2;159;89;55m \033[48;2;185;115;81m \033[48;2;200;130;96m \033[48;2;217;143;111m \033[48;2;212;141;110m \033[48;2;178;106;77m \033[48;2;178;107;78m \033[48;2;147;76;47m \033[m");
$display("\033[48;2;1;1;6m \033[48;2;0;0;5m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[48;2;5;6;9m \033[48;2;26;27;31m \033[48;2;24;27;32m \033[48;2;24;27;31m \033[48;2;20;23;30m \033[48;2;19;22;29m \033[48;2;19;22;31m \033[48;2;22;21;29m \033[48;2;10;9;15m \033[48;2;7;6;12m \033[48;2;5;4;9m \033[48;2;2;2;4m \033[48;2;2;2;4m \033[48;2;4;1;5m \033[48;2;4;2;5m \033[48;2;5;3;6m \033[48;2;10;5;12m \033[48;2;11;6;13m \033[48;2;10;5;12m \033[48;2;11;6;13m \033[48;2;12;7;14m \033[48;2;12;7;14m \033[48;2;13;8;15m \033[48;2;13;8;15m \033[48;2;13;8;15m \033[48;2;11;8;15m \033[48;2;15;10;14m \033[48;2;26;14;12m \033[48;2;98;72;65m \033[48;2;133;93;77m \033[48;2;151;109;85m \033[48;2;153;104;76m \033[48;2;157;103;73m \033[48;2;161;104;74m \033[48;2;161;102;70m \033[48;2;201;145;112m \033[48;2;227;172;138m \033[48;2;227;173;140m \033[48;2;229;171;138m \033[48;2;214;156;124m \033[48;2;209;145;118m \033[48;2;208;143;117m \033[48;2;211;145;121m \033[48;2;213;147;125m \033[48;2;208;142;122m \033[48;2;204;143;124m \033[48;2;195;136;121m \033[48;2;197;136;118m \033[48;2;202;141;123m \033[48;2;222;161;142m \033[48;2;244;183;162m \033[48;2;236;178;157m \033[48;2;231;176;155m \033[48;2;230;177;153m \033[48;2;248;193;170m \033[48;2;254;199;174m \033[48;2;252;199;173m \033[48;2;237;181;154m \033[48;2;200;143;116m \033[48;2;236;180;150m \033[48;2;226;170;143m \033[48;2;152;102;81m \033[48;2;81;48;29m \033[48;2;69;53;44m \033[48;2;62;57;57m \033[48;2;70;67;62m \033[48;2;71;67;64m \033[48;2;70;69;65m \033[48;2;70;69;66m \033[48;2;70;68;67m \033[48;2;70;66;67m \033[48;2;69;64;61m \033[48;2;64;56;52m \033[48;2;57;49;46m \033[48;2;60;52;49m \033[48;2;62;54;51m \033[48;2;64;56;54m \033[48;2;66;58;56m \033[48;2;67;58;59m \033[48;2;71;60;66m \033[48;2;69;62;66m \033[48;2;18;15;18m \033[48;2;15;15;17m \033[48;2;14;12;17m \033[48;2;6;4;9m \033[48;2;7;5;10m \033[48;2;12;3;10m \033[48;2;26;15;23m \033[48;2;42;23;34m \033[48;2;47;16;23m \033[48;2;176;139;119m \033[48;2;206;156;122m \033[48;2;162;84;52m \033[48;2;150;74;42m \033[48;2;154;84;50m \033[48;2;219;153;118m \033[48;2;201;134;100m \033[48;2;146;73;40m \033[48;2;145;72;38m \033[48;2;146;72;40m \033[48;2;207;134;101m \033[48;2;213;147;112m \033[48;2;140;75;41m \033[48;2;140;69;39m \033[48;2;139;66;38m \033[48;2;197;124;96m \033[m");
$display("\033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;2m \033[48;2;0;0;4m \033[48;2;22;23;28m \033[48;2;26;26;35m \033[48;2;33;36;45m \033[48;2;22;25;32m \033[48;2;20;22;30m \033[48;2;20;23;28m \033[48;2;10;14;18m \033[48;2;13;12;20m \033[48;2;9;8;14m \033[48;2;5;4;9m \033[48;2;1;0;5m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;1;1;1m \033[48;2;1;1;1m \033[48;2;1;1;1m \033[48;2;5;3;6m \033[48;2;6;4;9m \033[48;2;7;5;10m \033[48;2;7;4;11m \033[48;2;9;6;13m \033[48;2;9;6;13m \033[48;2;9;6;13m \033[48;2;9;6;13m \033[48;2;9;6;13m \033[48;2;14;11;18m \033[48;2;16;15;20m \033[48;2;100;88;88m \033[48;2;111;87;75m \033[48;2;120;79;62m \033[48;2;127;81;63m \033[48;2;150;99;80m \033[48;2;152;100;77m \033[48;2;155;101;77m \033[48;2;159;103;76m \033[48;2;178;119;90m \033[48;2;213;155;125m \033[48;2;230;177;143m \033[48;2;228;179;140m \033[48;2;231;173;138m \033[48;2;231;166;136m \033[48;2;223;161;132m \033[48;2;222;162;133m \033[48;2;223;160;132m \033[48;2;221;158;133m \033[48;2;221;160;137m \033[48;2;226;163;142m \033[48;2;226;174;152m \033[48;2;232;177;156m \033[48;2;235;177;157m \033[48;2;237;176;157m \033[48;2;236;175;156m \033[48;2;237;181;157m \033[48;2;247;193;167m \033[48;2;245;192;165m \033[48;2;244;192;164m \033[48;2;223;168;142m \033[48;2;190;134;107m \033[48;2;222;166;139m \033[48;2;194;136;113m \033[48;2;135;78;60m \033[48;2;83;39;26m \033[48;2;74;47;40m \033[48;2;65;54;51m \033[48;2;59;56;53m \033[48;2;60;59;55m \033[48;2;66;65;61m \033[48;2;73;70;65m \033[48;2;74;70;65m \033[48;2;75;70;64m \033[48;2;74;70;66m \033[48;2;76;71;68m \033[48;2;74;65;63m \033[48;2;62;54;52m \033[48;2;59;49;47m \033[48;2;61;53;50m \033[48;2;64;56;53m \033[48;2;64;58;54m \033[48;2;65;60;57m \033[48;2;65;59;61m \033[48;2;67;63;64m \033[48;2;43;41;45m \033[48;2;14;11;15m \033[48;2;17;15;18m \033[48;2;5;3;6m \033[48;2;5;3;6m \033[48;2;4;2;5m \033[48;2;13;7;12m \033[48;2;37;18;29m \033[48;2;53;21;26m \033[48;2;87;49;34m \033[48;2;189;134;108m \033[48;2;196;119;92m \033[48;2;136;60;31m \033[48;2;161;90;60m \033[48;2;198;131;99m \033[48;2;171;102;71m \033[48;2;133;59;28m \033[48;2;134;57;27m \033[48;2;137;61;31m \033[48;2;194;123;92m \033[48;2;192;127;94m \033[48;2;119;51;21m \033[48;2;120;51;22m \033[48;2;120;49;22m \033[48;2;146;78;47m \033[m");
$display("\033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;2m \033[48;2;12;11;15m \033[48;2;36;37;42m \033[48;2;38;38;46m \033[48;2;33;36;45m \033[48;2;22;25;32m \033[48;2;21;24;31m \033[48;2;6;9;14m \033[48;2;15;17;23m \033[48;2;6;6;13m \033[48;2;5;4;10m \033[48;2;1;0;6m \033[48;2;0;0;4m \033[48;2;0;0;2m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;2;0;3m \033[48;2;2;0;5m \033[48;2;3;1;6m \033[48;2;3;0;7m \033[48;2;9;0;11m \033[48;2;10;2;13m \033[48;2;10;2;13m \033[48;2;8;0;11m \033[48;2;25;16;28m \033[48;2;23;18;33m \033[48;2;16;15;29m \033[48;2;120;112;120m \033[48;2;100;78;80m \033[48;2;110;73;63m \033[48;2;115;67;57m \033[48;2;120;63;50m \033[48;2;138;84;63m \033[48;2;149;101;75m \033[48;2;156;102;78m \033[48;2;175;117;93m \033[48;2;208;152;125m \033[48;2;236;184;153m \033[48;2;248;198;166m \033[48;2;250;199;168m \033[48;2;245;195;165m \033[48;2;242;192;165m \033[48;2;244;194;168m \033[48;2;244;197;170m \033[48;2;250;204;179m \033[48;2;255;209;186m \033[48;2;255;210;188m \033[48;2;251;207;183m \033[48;2;248;201;179m \033[48;2;247;200;177m \033[48;2;249;201;179m \033[48;2;249;203;179m \033[48;2;249;203;177m \033[48;2;249;202;174m \033[48;2;240;190;163m \033[48;2;218;167;138m \033[48;2;188;129;108m \033[48;2;205;152;128m \033[48;2;149;104;80m \033[48;2;101;61;43m \033[48;2;61;28;14m \033[48;2;70;46;36m \033[48;2;64;49;43m \033[48;2;57;50;47m \033[48;2;65;62;57m \033[48;2;72;71;66m \033[48;2;81;80;75m \033[48;2;92;89;82m \033[48;2;90;85;77m \033[48;2;82;79;72m \033[48;2;73;69;66m \033[48;2;63;58;55m \033[48;2;62;54;51m \033[48;2;60;52;50m \033[48;2;59;48;46m \033[48;2;58;50;47m \033[48;2;63;55;52m \033[48;2;62;57;53m \033[48;2;64;59;56m \033[48;2;67;61;63m \033[48;2;66;62;63m \033[48;2;63;61;64m \033[48;2;10;8;11m \033[48;2;17;15;18m \033[48;2;12;10;13m \033[48;2;2;0;3m \033[48;2;2;0;3m \033[48;2;10;6;9m \033[48;2;26;12;15m \033[48;2;43;24;22m \033[48;2;50;18;13m \033[48;2;107;55;37m \033[48;2;127;55;31m \033[48;2;124;52;28m \033[48;2;123;53;28m \033[48;2;126;56;31m \033[48;2;125;54;30m \033[48;2;124;50;26m \033[48;2;123;47;25m \033[48;2;120;45;21m \033[48;2;120;51;26m \033[48;2;117;47;20m \033[48;2;116;44;20m \033[48;2;118;46;23m \033[48;2;120;45;23m \033[48;2;117;47;22m \033[m");
$display("\033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;1m \033[48;2;49;48;54m \033[48;2;34;34;42m \033[48;2;48;48;59m \033[48;2;31;34;43m \033[48;2;13;16;23m \033[48;2;11;14;21m \033[48;2;4;7;12m \033[48;2;1;3;8m \033[48;2;2;1;6m \033[48;2;0;0;4m \033[48;2;0;0;4m \033[48;2;0;0;4m \033[48;2;1;1;4m \033[48;2;1;0;5m \033[48;2;1;0;5m \033[48;2;1;0;6m \033[48;2;1;0;6m \033[48;2;3;0;6m \033[48;2;1;0;5m \033[48;2;1;1;7m \033[48;2;1;1;9m \033[48;2;2;1;9m \033[48;2;12;11;19m \033[48;2;23;21;30m \033[48;2;27;24;35m \033[48;2;23;18;32m \033[48;2;16;14;31m \033[48;2;24;22;41m \033[48;2;114;109;123m \033[48;2;105;91;99m \033[48;2;90;53;54m \033[48;2;106;56;43m \033[48;2;111;53;32m \033[48;2;107;51;28m \033[48;2;112;61;34m \033[48;2;132;80;56m \033[48;2;148;96;69m \033[48;2;163;113;85m \033[48;2;194;145;115m \033[48;2;227;180;150m \033[48;2;239;193;165m \033[48;2;246;201;172m \033[48;2;246;202;175m \033[48;2;243;201;173m \033[48;2;243;203;172m \033[48;2;244;199;172m \033[48;2;238;196;170m \033[48;2;247;209;183m \033[48;2;252;217;189m \033[48;2;249;212;185m \033[48;2;246;206;180m \033[48;2;248;205;180m \033[48;2;247;205;177m \033[48;2;247;203;174m \033[48;2;235;189;162m \033[48;2;202;153;126m \033[48;2;171;121;89m \033[48;2;175;122;101m \033[48;2;122;76;68m \033[48;2;71;38;33m \033[48;2;61;43;36m \033[48;2;46;34;32m \033[48;2;63;55;50m \033[48;2;53;47;43m \033[48;2;64;59;56m \033[48;2;67;64;63m \033[48;2;68;63;60m \033[48;2;75;70;66m \033[48;2;81;77;72m \033[48;2;80;75;71m \033[48;2;65;60;56m \033[48;2;53;48;44m \033[48;2;38;33;29m \033[48;2;23;18;15m \033[48;2;16;11;8m \033[48;2;56;48;46m \033[48;2;55;47;44m \033[48;2;63;55;52m \033[48;2;64;57;51m \033[48;2;65;58;52m \033[48;2;67;62;58m \033[48;2;68;62;61m \033[48;2;66;62;63m \033[48;2;45;41;42m \033[48;2;18;13;17m \033[48;2;17;12;16m \033[48;2;6;1;5m \033[48;2;4;0;3m \033[48;2;6;1;6m \033[48;2;18;12;15m \033[48;2;33;26;25m \033[48;2;42;24;18m \033[48;2;92;55;45m \033[48;2;122;63;50m \033[48;2;139;80;67m \033[48;2;137;78;65m \033[48;2;143;84;71m \033[48;2;111;52;39m \033[48;2;111;47;37m \033[48;2;110;46;36m \033[48;2;108;45;34m \033[48;2;102;38;28m \033[48;2;112;47;37m \033[48;2;133;68;56m \033[48;2;110;45;32m \033[48;2;110;45;32m \033[48;2;111;44;33m \033[m");
$display("\033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;17;17;18m \033[48;2;74;73;80m \033[48;2;35;35;45m \033[48;2;61;61;72m \033[48;2;25;29;38m \033[48;2;5;8;15m \033[48;2;3;6;13m \033[48;2;10;13;18m \033[48;2;0;0;5m \033[48;2;0;0;5m \033[48;2;0;0;4m \033[48;2;0;0;4m \033[48;2;0;0;4m \033[48;2;3;2;7m \033[48;2;10;9;14m \033[48;2;19;19;24m \033[48;2;25;24;32m \033[48;2;29;28;36m \033[48;2;30;28;39m \033[48;2;31;31;40m \033[48;2;27;28;40m \033[48;2;26;28;40m \033[48;2;25;25;37m \033[48;2;23;23;35m \033[48;2;24;21;35m \033[48;2;24;22;36m \033[48;2;20;17;33m \033[48;2;17;14;33m \033[48;2;33;30;47m \033[48;2;112;108;123m \033[48;2;114;108;121m \033[48;2;118;94;96m \033[48;2;75;41;35m \033[48;2;93;47;25m \033[48;2;102;50;19m \033[48;2;108;53;27m \033[48;2;102;50;26m \033[48;2;100;49;22m \033[48;2;117;68;40m \033[48;2;130;80;51m \033[48;2;149;100;70m \033[48;2;185;135;108m \033[48;2;201;153;126m \033[48;2;220;173;147m \033[48;2;234;189;163m \033[48;2;238;194;167m \033[48;2;239;193;164m \033[48;2;220;174;146m \033[48;2;209;167;135m \033[48;2;223;185;151m \033[48;2;230;189;159m \033[48;2;238;194;167m \033[48;2;235;188;165m \033[48;2;232;183;160m \033[48;2;220;174;147m \033[48;2;188;141;113m \033[48;2;140;93;67m \033[48;2;116;68;47m \033[48;2;83;42;32m \033[48;2;70;41;41m \033[48;2;38;28;25m \033[48;2;51;51;45m \033[48;2;42;43;46m \033[48;2;40;40;44m \033[48;2;58;56;59m \033[48;2;55;53;54m \033[48;2;55;51;52m \033[48;2;55;48;48m \033[48;2;57;51;51m \033[48;2;62;56;56m \033[48;2;51;45;45m \033[48;2;36;30;30m \033[48;2;20;14;14m \033[48;2;7;1;1m \033[48;2;6;0;0m \033[48;2;7;1;1m \033[48;2;57;49;47m \033[48;2;54;47;43m \033[48;2;60;52;49m \033[48;2;63;56;49m \033[48;2;64;57;51m \033[48;2;66;61;55m \033[48;2;67;62;58m \033[48;2;67;63;61m \033[48;2;66;62;61m \033[48;2;19;14;19m \033[48;2;18;13;17m \033[48;2;11;6;10m \033[48;2;6;1;5m \033[48;2;5;0;3m \033[48;2;12;6;8m \033[48;2;29;23;20m \033[48;2;36;22;19m \033[48;2;38;19;17m \033[48;2;33;7;2m \033[48;2;34;7;3m \033[48;2;35;7;2m \033[48;2;34;6;1m \033[48;2;33;6;2m \033[48;2;33;8;7m \033[48;2;40;13;12m \033[48;2;35;10;8m \033[48;2;26;0;0m \033[48;2;21;0;0m \033[48;2;24;1;2m \033[48;2;26;4;3m \033[48;2;26;4;3m \033[48;2;25;3;1m \033[m");
$display("\033[48;2;0;0;0m \033[48;2;0;1;0m \033[48;2;53;57;60m \033[48;2;66;70;75m \033[48;2;41;44;52m \033[48;2;60;62;74m \033[48;2;14;15;21m \033[48;2;6;6;11m \033[48;2;0;0;4m \033[48;2;6;6;12m \033[48;2;0;0;4m \033[48;2;10;9;13m \033[48;2;18;16;22m \033[48;2;21;19;29m \033[48;2;23;20;34m \033[48;2;19;21;33m \033[48;2;19;21;33m \033[48;2;20;22;34m \033[48;2;21;23;35m \033[48;2;23;25;37m \033[48;2;27;29;41m \033[48;2;28;30;42m \033[48;2;30;32;44m \033[48;2;33;35;47m \033[48;2;35;37;49m \033[48;2;36;38;50m \033[48;2;37;39;51m \033[48;2;35;37;49m \033[48;2;26;28;40m \033[48;2;17;19;30m \033[48;2;20;23;34m \033[48;2;103;105;116m \033[48;2;110;113;124m \033[48;2;114;112;125m \033[48;2;116;106;116m \033[48;2;83;62;63m \033[48;2;59;27;15m \033[48;2;86;49;27m \033[48;2;99;54;28m \033[48;2;100;52;22m \033[48;2;101;51;25m \033[48;2;98;48;28m \033[48;2;97;44;21m \033[48;2;94;42;20m \033[48;2;95;46;25m \033[48;2;95;47;26m \033[48;2;104;58;39m \033[48;2;130;84;65m \033[48;2;155;109;92m \033[48;2;157;111;93m \033[48;2;140;95;76m \033[48;2;137;94;76m \033[48;2;139;93;77m \033[48;2;138;89;74m \033[48;2;139;89;73m \033[48;2;127;76;62m \033[48;2;106;56;46m \033[48;2;108;58;48m \033[48;2;104;58;42m \033[48;2;94;51;44m \033[48;2;35;2;5m \033[48;2;52;34;49m \033[48;2;83;81;94m \033[48;2;49;51;61m \033[48;2;48;46;60m \033[48;2;42;42;50m \033[48;2;51;50;56m \033[48;2;48;47;51m \033[48;2;45;43;46m \033[48;2;38;38;39m \033[48;2;19;20;20m \033[48;2;6;6;7m \033[48;2;4;4;6m \033[48;2;2;2;3m \033[48;2;1;1;3m \033[48;2;3;3;5m \033[48;2;12;10;13m \033[48;2;11;8;12m \033[48;2;25;19;26m \033[48;2;35;29;33m \033[48;2;45;39;39m \033[48;2;62;54;51m \033[48;2;64;57;54m \033[48;2;66;58;55m \033[48;2;69;61;58m \033[48;2;71;63;61m \033[48;2;71;63;61m \033[48;2;45;35;38m \033[48;2;21;12;15m \033[48;2;17;7;11m \033[48;2;9;0;3m \033[48;2;7;1;3m \033[48;2;4;0;3m \033[48;2;21;15;15m \033[48;2;34;21;20m \033[48;2;39;16;17m \033[48;2;45;16;19m \033[48;2;51;20;16m \033[48;2;59;28;23m \033[48;2;59;30;10m \033[48;2;61;29;20m \033[48;2;44;16;3m \033[48;2;87;61;44m \033[48;2;77;49;35m \033[48;2;42;18;10m \033[48;2;35;22;11m \033[48;2;27;17;7m \033[48;2;22;11;3m \033[48;2;21;11;2m \033[48;2;20;10;2m \033[m");
$display("\033[48;2;0;0;2m \033[48;2;2;4;6m \033[48;2;32;36;39m \033[48;2;30;33;38m \033[48;2;31;34;39m \033[48;2;15;18;23m \033[48;2;1;2;5m \033[48;2;4;4;8m \033[48;2;6;7;11m \033[48;2;20;20;25m \033[48;2;21;22;26m \033[48;2;21;24;31m \033[48;2;20;23;30m \033[48;2;21;24;33m \033[48;2;20;23;32m \033[48;2;19;23;34m \033[48;2;19;23;34m \033[48;2;25;28;39m \033[48;2;27;31;42m \033[48;2;29;33;44m \033[48;2;30;35;46m \033[48;2;32;36;47m \033[48;2;33;37;48m \033[48;2;36;40;51m \033[48;2;38;42;53m \033[48;2;38;42;53m \033[48;2;40;44;55m \033[48;2;41;45;56m \033[48;2;41;45;56m \033[48;2;33;37;48m \033[48;2;22;26;37m \033[48;2;73;77;88m \033[48;2;109;113;124m \033[48;2;110;114;125m \033[48;2;113;113;123m \033[48;2;120;114;117m \033[48;2;96;85;80m \033[48;2;80;61;48m \033[48;2;58;23;5m \033[48;2;94;52;29m \033[48;2;103;54;26m \033[48;2;105;56;26m \033[48;2;107;57;32m \033[48;2;105;57;35m \033[48;2;104;58;40m \033[48;2;88;45;31m \033[48;2;83;43;33m \033[48;2;78;42;30m \033[48;2;78;40;29m \033[48;2;78;40;29m \033[48;2;79;42;31m \033[48;2;75;42;31m \033[48;2;87;48;40m \033[48;2;101;54;48m \033[48;2;109;57;53m \033[48;2;110;55;49m \033[48;2;110;56;46m \033[48;2;110;53;46m \033[48;2;94;49;37m \033[48;2;43;9;4m \033[48;2;22;0;8m \033[48;2;155;138;163m \033[48;2;102;96;120m \033[48;2;30;30;42m \033[48;2;28;28;38m \033[48;2;38;38;48m \033[48;2;28;28;36m \033[48;2;24;24;29m \033[48;2;4;2;8m \033[48;2;1;1;3m \033[48;2;0;1;2m \033[48;2;2;2;4m \033[48;2;1;1;3m \033[48;2;5;4;6m \033[48;2;8;7;12m \033[48;2;12;11;16m \033[48;2;16;15;19m \033[48;2;18;16;21m \033[48;2;16;14;19m \033[48;2;21;16;20m \033[48;2;29;25;24m \033[48;2;39;34;31m \033[48;2;55;50;46m \033[48;2;64;56;53m \033[48;2;68;60;57m \033[48;2;71;63;61m \033[48;2;71;63;61m \033[48;2;63;54;57m \033[48;2;21;12;15m \033[48;2;17;8;11m \033[48;2;10;1;4m \033[48;2;6;0;2m \033[48;2;4;0;3m \033[48;2;19;13;13m \033[48;2;31;17;17m \033[48;2;40;17;20m \033[48;2;143;108;40m \033[48;2;255;217;64m \033[48;2;237;179;26m \033[48;2;228;167;25m \033[48;2;231;163;21m \033[48;2;165;92;1m \033[48;2;149;84;28m \033[48;2;131;71;28m \033[48;2;171;112;47m \033[48;2;119;69;23m \033[48;2;39;14;1m \033[48;2;22;11;7m \033[48;2;19;13;4m \033[48;2;17;14;2m \033[m");
$display("\033[48;2;40;41;46m \033[48;2;38;38;46m \033[48;2;30;34;40m \033[48;2;23;27;33m \033[48;2;22;27;32m \033[48;2;22;27;31m \033[48;2;22;25;30m \033[48;2;22;25;30m \033[48;2;23;26;32m \033[48;2;24;27;32m \033[48;2;25;28;35m \033[48;2;23;27;36m \033[48;2;22;26;35m \033[48;2;22;26;35m \033[48;2;22;26;35m \033[48;2;19;22;31m \033[48;2;30;33;42m \033[48;2;30;32;44m \033[48;2;30;32;44m \033[48;2;31;33;46m \033[48;2;32;36;47m \033[48;2;37;41;52m \033[48;2;37;41;52m \033[48;2;40;44;55m \033[48;2;39;43;54m \033[48;2;39;43;54m \033[48;2;38;42;54m \033[48;2;37;41;53m \033[48;2;35;38;53m \033[48;2;38;41;58m \033[48;2;39;42;58m \033[48;2;41;44;60m \033[48;2;89;92;108m \033[48;2;114;114;132m \033[48;2;114;113;128m \033[48;2;115;113;125m \033[48;2;114;113;119m \033[48;2;97;92;94m \033[48;2;87;74;68m \033[48;2;74;52;38m \033[48;2;53;20;0m \033[48;2;83;46;20m \033[48;2;103;57;34m \033[48;2;105;58;38m \033[48;2;107;56;35m \033[48;2;107;56;34m \033[48;2;108;56;34m \033[48;2;107;55;34m \033[48;2;112;60;39m \033[48;2;114;59;39m \033[48;2;117;59;41m \033[48;2;118;55;38m \033[48;2;115;51;36m \033[48;2;122;58;44m \033[48;2;125;59;47m \033[48;2;125;59;47m \033[48;2;116;53;44m \033[48;2;113;54;48m \033[48;2;65;17;13m \033[48;2;27;1;1m \033[48;2;85;68;94m \033[48;2;182;166;203m \033[48;2;52;42;71m \033[48;2;31;30;43m \033[48;2;30;30;38m \033[48;2;27;25;38m \033[48;2;28;26;36m \033[48;2;29;28;36m \033[48;2;32;31;39m \033[48;2;24;23;29m \033[48;2;1;1;7m \033[48;2;47;46;52m \033[48;2;13;12;18m \033[48;2;13;12;18m \033[48;2;12;10;19m \033[48;2;13;11;22m \033[48;2;17;16;24m \033[48;2;17;16;24m \033[48;2;15;13;18m \033[48;2;17;15;20m \033[48;2;29;25;29m \033[48;2;38;33;30m \033[48;2;48;41;36m \033[48;2;59;52;46m \033[48;2;65;59;53m \033[48;2;69;61;58m \033[48;2;72;64;61m \033[48;2;75;66;68m \033[48;2;37;27;29m \033[48;2;18;11;13m \033[48;2;10;3;5m \033[48;2;5;1;1m \033[48;2;4;0;1m \033[48;2;8;3;3m \033[48;2;28;15;15m \033[48;2;40;20;21m \033[48;2;63;17;10m \033[48;2;165;84;14m \033[48;2;168;64;3m \033[48;2;169;66;6m \033[48;2;168;58;6m \033[48;2;155;50;4m \033[48;2;150;76;36m \033[48;2;122;54;20m \033[48;2;127;55;9m \033[48;2;88;36;4m \033[48;2;32;14;3m \033[48;2;21;13;10m \033[48;2;22;14;3m \033[48;2;18;15;6m \033[m");
$display("\033[48;2;41;41;48m \033[48;2;37;40;47m \033[48;2;30;35;41m \033[48;2;23;28;34m \033[48;2;24;29;35m \033[48;2;23;28;34m \033[48;2;23;26;33m \033[48;2;23;26;33m \033[48;2;24;27;34m \033[48;2;24;27;34m \033[48;2;25;28;35m \033[48;2;24;28;37m \033[48;2;24;28;37m \033[48;2;24;28;37m \033[48;2;23;27;36m \033[48;2;22;26;35m \033[48;2;17;21;31m \033[48;2;2;6;16m \033[48;2;23;27;38m \033[48;2;31;35;47m \033[48;2;38;42;53m \033[48;2;38;42;53m \033[48;2;35;39;50m \033[48;2;34;38;49m \033[48;2;32;36;47m \033[48;2;32;36;47m \033[48;2;31;35;47m \033[48;2;33;37;51m \033[48;2;36;39;54m \033[48;2;39;42;61m \033[48;2;43;46;65m \033[48;2;43;46;65m \033[48;2;70;73;92m \033[48;2;105;106;126m \033[48;2;110;111;129m \033[48;2;114;116;131m \033[48;2;112;114;127m \033[48;2;107;110;122m \033[48;2;88;88;95m \033[48;2;81;75;85m \033[48;2;82;67;68m \033[48;2;78;56;43m \033[48;2;66;33;14m \033[48;2;92;52;32m \033[48;2;99;55;32m \033[48;2;104;54;28m \033[48;2;107;54;25m \033[48;2;115;59;29m \033[48;2;127;68;40m \033[48;2;135;71;44m \033[48;2;138;72;46m \033[48;2;138;74;47m \033[48;2;129;65;39m \033[48;2;125;60;38m \033[48;2;125;60;41m \033[48;2;125;58;43m \033[48;2;118;55;43m \033[48;2;98;46;40m \033[48;2;36;2;11m \033[48;2;173;149;180m \033[48;2;197;183;233m \033[48;2;149;137;182m \033[48;2;38;30;65m \033[48;2;34;31;51m \033[48;2;31;30;44m \033[48;2;28;26;39m \033[48;2;24;22;35m \033[48;2;25;23;34m \033[48;2;22;20;31m \033[48;2;27;25;36m \033[48;2;31;29;40m \033[48;2;25;24;32m \033[48;2;17;16;23m \033[48;2;13;11;20m \033[48;2;12;10;21m \033[48;2;13;11;22m \033[48;2;14;13;20m \033[48;2;14;13;20m \033[48;2;15;13;17m \033[48;2;12;9;16m \033[48;2;28;23;29m \033[48;2;37;32;32m \033[48;2;45;40;34m \033[48;2;53;46;38m \033[48;2;59;52;46m \033[48;2;67;60;56m \033[48;2;71;63;60m \033[48;2;71;63;61m \033[48;2;66;57;58m \033[48;2;21;15;16m \033[48;2;18;13;15m \033[48;2;2;0;0m \033[48;2;1;0;0m \033[48;2;8;4;3m \033[48;2;24;15;13m \033[48;2;37;20;20m \033[48;2;55;21;15m \033[48;2;201;165;70m \033[48;2;226;200;22m \033[48;2;233;210;38m \033[48;2;238;216;33m \033[48;2;229;198;58m \033[48;2;129;69;6m \033[48;2;197;105;68m \033[48;2;143;51;23m \033[48;2;70;33;9m \033[48;2;32;17;7m \033[48;2;20;15;9m \033[48;2;19;16;6m \033[48;2;20;17;9m \033[m");
$display("\033[48;2;27;27;34m \033[48;2;27;27;35m \033[48;2;26;29;36m \033[48;2;24;27;34m \033[48;2;25;28;35m \033[48;2;25;28;35m \033[48;2;27;30;39m \033[48;2;27;30;39m \033[48;2;27;30;39m \033[48;2;27;30;39m \033[48;2;27;30;39m \033[48;2;26;30;39m \033[48;2;26;30;39m \033[48;2;26;30;39m \033[48;2;26;30;39m \033[48;2;32;35;43m \033[48;2;26;29;38m \033[48;2;27;29;41m \033[48;2;34;36;48m \033[48;2;31;33;45m \033[48;2;32;36;47m \033[48;2;32;36;47m \033[48;2;32;36;47m \033[48;2;32;36;47m \033[48;2;33;37;48m \033[48;2;33;37;48m \033[48;2;34;38;50m \033[48;2;36;40;53m \033[48;2;39;43;59m \033[48;2;45;47;68m \033[48;2;48;50;71m \033[48;2;42;44;65m \033[48;2;54;57;77m \033[48;2;88;92;110m \033[48;2;110;113;132m \033[48;2;114;117;136m \033[48;2;117;120;139m \033[48;2;119;122;141m \033[48;2;118;118;140m \033[48;2;93;96;108m \033[48;2;94;91;96m \033[48;2;101;86;85m \033[48;2;108;83;82m \033[48;2;113;81;75m \033[48;2;101;59;48m \033[48;2;87;36;19m \033[48;2;103;46;23m \033[48;2;117;63;37m \033[48;2;121;62;39m \033[48;2;125;64;41m \033[48;2;126;62;39m \033[48;2;125;60;40m \033[48;2;126;61;43m \033[48;2;126;60;43m \033[48;2;136;70;56m \033[48;2;158;95;83m \033[48;2;157;101;100m \033[48;2;146;104;125m \033[48;2;211;194;233m \033[48;2;202;196;244m \033[48;2;158;150;202m \033[48;2;133;127;167m \033[48;2;35;30;60m \033[48;2;45;42;60m \033[48;2;41;39;51m \033[48;2;34;33;47m \033[48;2;29;27;41m \033[48;2;26;24;37m \033[48;2;27;25;38m \033[48;2;27;25;38m \033[48;2;29;27;40m \033[48;2;29;27;38m \033[48;2;10;8;19m \033[48;2;12;11;20m \033[48;2;12;10;21m \033[48;2;13;11;22m \033[48;2;13;12;20m \033[48;2;13;12;20m \033[48;2;13;10;17m \033[48;2;12;9;18m \033[48;2;14;9;16m \033[48;2;38;33;34m \033[48;2;47;42;37m \033[48;2;52;45;39m \033[48;2;60;53;47m \033[48;2;68;60;57m \033[48;2;70;62;59m \033[48;2;73;64;65m \033[48;2;79;70;71m \033[48;2;20;14;16m \033[48;2;20;15;16m \033[48;2;3;0;1m \033[48;2;1;1;1m \033[48;2;168;122;172m \033[48;2;169;121;172m \033[48;2;171;120;171m \033[48;2;172;119;170m \033[48;2;166;112;155m \033[48;2;156;100;84m \033[48;2;116;57;29m \033[48;2;86;27;5m \033[48;2;133;69;43m \033[48;2;116;65;42m \033[48;2;67;13;2m \033[48;2;50;15;0m \033[48;2;35;16;0m \033[48;2;29;19;8m \033[48;2;18;15;10m \033[48;2;16;16;9m \033[48;2;20;16;9m \033[m");
$display("\033[48;2;30;29;36m \033[48;2;30;28;36m \033[48;2;30;30;38m \033[48;2;30;32;40m \033[48;2;32;35;42m \033[48;2;33;36;43m \033[48;2;33;36;43m \033[48;2;33;36;43m \033[48;2;32;35;43m \033[48;2;35;38;45m \033[48;2;31;34;41m \033[48;2;173;119;170m \033[48;2;172;120;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;167;122;173m \033[48;2;165;123;173m \033[48;2;163;124;174m \033[48;2;162;125;175m \033[48;2;160;126;176m \033[48;2;158;127;176m \033[48;2;156;128;177m \033[48;2;154;129;178m \033[48;2;35;39;50m \033[48;2;34;38;49m \033[48;2;36;40;52m \033[48;2;39;42;56m \033[48;2;39;42;59m \033[48;2;44;47;66m \033[48;2;48;51;73m \033[48;2;48;51;74m \033[48;2;29;31;55m \033[48;2;58;60;85m \033[48;2;67;69;94m \033[48;2;129;138;182m \033[48;2;129;142;188m \033[48;2;128;143;189m \033[48;2;126;144;189m \033[48;2;124;145;190m \033[48;2;123;145;191m \033[48;2;121;146;191m \033[48;2;133;121;129m \033[48;2;121;107;115m \033[48;2;112;95;104m \033[48;2;115;93;98m \033[48;2;120;93;88m \033[48;2;102;69;58m \033[48;2;71;36;18m \033[48;2;80;42;24m \033[48;2;89;45;24m \033[48;2;103;54;32m \033[48;2;116;67;53m \033[48;2;109;153;196m \033[48;2;108;153;196m \033[48;2;108;153;196m \033[48;2;108;153;196m \033[48;2;109;153;196m \033[48;2;109;153;196m \033[48;2;109;152;196m \033[48;2;110;152;196m \033[48;2;111;152;195m \033[48;2;112;151;195m \033[48;2;113;151;195m \033[48;2;46;46;64m \033[48;2;53;55;69m \033[48;2;56;54;68m \033[48;2;43;41;55m \033[48;2;41;40;53m \033[48;2;41;39;53m \033[48;2;41;37;51m \033[48;2;39;37;48m \033[48;2;126;144;189m \033[48;2;127;143;189m \033[48;2;129;142;188m \033[48;2;131;141;187m \033[48;2;133;140;186m \033[48;2;135;139;186m \033[48;2;137;138;185m \033[48;2;138;137;184m \033[48;2;140;136;183m \033[48;2;142;135;183m \033[48;2;144;134;182m \033[48;2;39;34;37m \033[48;2;46;38;38m \033[48;2;61;53;51m \033[48;2;66;59;56m \033[48;2;68;61;58m \033[48;2;65;61;60m \033[48;2;67;63;61m \033[48;2;46;42;44m \033[48;2;22;18;19m \033[48;2;8;6;7m \033[48;2;1;1;1m \033[48;2;167;122;173m \033[48;2;168;121;172m \033[48;2;170;120;171m \033[48;2;172;120;171m \033[48;2;90;60;82m \033[48;2;33;18;14m \033[48;2;35;19;15m \033[48;2;45;28;22m \033[48;2;47;27;24m \033[48;2;54;34;33m \033[48;2;33;18;19m \033[48;2;27;18;17m \033[48;2;25;17;14m \033[48;2;24;17;13m \033[48;2;19;14;10m \033[48;2;18;13;9m \033[48;2;32;28;25m \033[m");
$display("\033[48;2;34;30;39m \033[48;2;36;33;42m \033[48;2;35;34;42m \033[48;2;36;35;43m \033[48;2;36;36;45m \033[48;2;37;37;45m \033[48;2;36;39;44m \033[48;2;36;39;44m \033[48;2;36;39;44m \033[48;2;35;38;43m \033[48;2;34;37;42m \033[48;2;173;119;170m \033[48;2;171;120;171m \033[48;2;169;121;172m \033[48;2;168;122;172m \033[48;2;166;123;173m \033[48;2;164;123;174m \033[48;2;162;124;175m \033[48;2;161;125;175m \033[48;2;159;126;176m \033[48;2;157;127;177m \033[48;2;155;128;178m \033[48;2;153;129;178m \033[48;2;151;130;179m \033[48;2;149;131;180m \033[48;2;69;66;91m \033[48;2;43;46;63m \033[48;2;45;48;67m \033[48;2;50;51;72m \033[48;2;50;56;78m \033[48;2;51;55;80m \033[48;2;45;49;75m \033[48;2;42;46;72m \033[48;2;69;73;102m \033[48;2;130;142;188m \033[48;2;128;143;189m \033[48;2;126;144;189m \033[48;2;124;145;190m \033[48;2;122;146;191m \033[48;2;121;146;191m \033[48;2;119;147;192m \033[48;2;134;144;176m \033[48;2;148;141;164m \033[48;2;146;142;166m \033[48;2;144;142;164m \033[48;2;143;136;156m \033[48;2;149;136;155m \033[48;2;137;118;135m \033[48;2;122;102;115m \033[48;2;78;45;55m \033[48;2;107;154;197m \033[48;2;106;154;197m \033[48;2;106;154;197m \033[48;2;105;155;198m \033[48;2;105;155;198m \033[48;2;105;155;198m \033[48;2;106;154;197m \033[48;2;106;154;197m \033[48;2;107;154;197m \033[48;2;107;153;197m \033[48;2;108;153;196m \033[48;2;109;152;196m \033[48;2;110;152;196m \033[48;2;250;248;254m \033[48;2;254;254;254m \033[48;2;254;253;255m \033[48;2;245;244;250m \033[48;2;170;169;175m \033[48;2;75;74;79m \033[48;2;121;146;191m \033[48;2;122;146;191m \033[48;2;124;145;190m \033[48;2;126;144;189m \033[48;2;128;143;189m \033[48;2;129;142;188m \033[48;2;131;141;187m \033[48;2;133;140;186m \033[48;2;135;139;186m \033[48;2;137;138;185m \033[48;2;139;137;184m \033[48;2;141;136;183m \033[48;2;143;135;182m \033[48;2;28;25;31m \033[48;2;34;29;33m \033[48;2;31;28;28m \033[48;2;34;30;31m \033[48;2;41;37;36m \033[48;2;52;51;49m \033[48;2;59;58;56m \033[48;2;60;58;58m \033[48;2;14;12;13m \033[48;2;11;10;11m \033[48;2;1;0;2m \033[48;2;166;123;173m \033[48;2;168;122;172m \033[48;2;169;121;172m \033[48;2;171;120;171m \033[48;2;28;18;17m \033[48;2;41;25;26m \033[48;2;45;27;27m \033[48;2;55;34;34m \033[48;2;58;40;38m \033[48;2;37;19;19m \033[48;2;19;5;7m \033[48;2;16;11;11m \033[48;2;20;14;14m \033[48;2;19;13;13m \033[48;2;18;14;13m \033[48;2;18;14;13m \033[48;2;29;25;24m \033[m");
$display("\033[48;2;37;35;40m \033[48;2;39;36;43m \033[48;2;39;38;44m \033[48;2;41;40;46m \033[48;2;41;42;47m \033[48;2;42;43;48m \033[48;2;39;42;47m \033[48;2;39;42;47m \033[48;2;38;41;46m \033[48;2;38;41;46m \033[48;2;37;40;44m \033[48;2;172;119;171m \033[48;2;171;120;171m \033[48;2;169;121;172m \033[48;2;167;122;173m \033[48;2;48;49;58m \033[48;2;39;43;52m \033[48;2;42;46;55m \033[48;2;43;47;56m \033[48;2;44;48;59m \033[48;2;45;49;61m \033[48;2;92;83;110m \033[48;2;152;130;179m \033[48;2;150;131;179m \033[48;2;148;132;180m \033[48;2;146;133;181m \033[48;2;46;49;68m \033[48;2;50;52;73m \033[48;2;53;55;76m \033[48;2;60;62;85m \033[48;2;56;59;82m \033[48;2;47;51;76m \033[48;2;46;50;75m \033[48;2;130;141;187m \033[48;2;128;142;188m \033[48;2;126;143;189m \033[48;2;125;144;190m \033[48;2;159;162;196m \033[48;2;121;146;191m \033[48;2;119;147;192m \033[48;2;118;148;193m \033[48;2;116;149;193m \033[48;2;214;215;245m \033[48;2;221;222;250m \033[48;2;228;228;253m \033[48;2;231;231;254m \033[48;2;233;233;254m \033[48;2;232;231;252m \033[48;2;218;206;229m \033[48;2;105;155;198m \033[48;2;104;155;198m \033[48;2;104;155;198m \033[48;2;103;156;199m \033[48;2;103;156;199m \033[48;2;157;123;157m \033[48;2;232;216;250m \033[48;2;208;206;242m \033[48;2;195;196;243m \033[48;2;188;189;233m \033[48;2;177;176;219m \033[48;2;159;152;191m \033[48;2;227;224;245m \033[48;2;253;253;255m \033[48;2;255;255;254m \033[48;2;252;252;250m \033[48;2;254;254;254m \033[48;2;254;254;254m \033[48;2;254;254;254m \033[48;2;120;150;194m \033[48;2;119;147;192m \033[48;2;121;146;191m \033[48;2;123;145;191m \033[48;2;124;144;190m \033[48;2;15;15;25m \033[48;2;11;11;24m \033[48;2;11;11;23m \033[48;2;9;11;22m \033[48;2;8;10;22m \033[48;2;7;9;21m \033[48;2;8;10;21m \033[48;2;13;12;20m \033[48;2;31;28;35m \033[48;2;35;33;38m \033[48;2;35;33;38m \033[48;2;37;32;38m \033[48;2;36;31;37m \033[48;2;35;28;35m \033[48;2;35;30;36m \033[48;2;32;27;33m \033[48;2;31;29;32m \033[48;2;26;25;27m \033[48;2;22;20;23m \033[48;2;2;1;4m \033[48;2;165;123;173m \033[48;2;167;122;173m \033[48;2;169;121;172m \033[48;2;170;120;171m \033[48;2;27;19;17m \033[48;2;37;27;25m \033[48;2;75;64;62m \033[48;2;74;57;57m \033[48;2;63;44;46m \033[48;2;45;30;33m \033[48;2;40;28;32m \033[48;2;31;21;26m \033[48;2;22;16;21m \033[48;2;17;11;12m \033[48;2;12;8;5m \033[48;2;10;6;4m \033[48;2;15;11;12m \033[m");
$display("\033[48;2;41;39;45m \033[48;2;43;40;47m \033[48;2;41;40;46m \033[48;2;42;41;47m \033[48;2;42;43;48m \033[48;2;43;44;49m \033[48;2;42;45;52m \033[48;2;41;44;51m \033[48;2;41;44;51m \033[48;2;40;43;50m \033[48;2;40;43;50m \033[48;2;172;119;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;167;122;173m \033[48;2;48;50;59m \033[48;2;42;46;55m \033[48;2;45;49;58m \033[48;2;45;49;59m \033[48;2;47;51;62m \033[48;2;49;52;67m \033[48;2;51;54;69m \033[48;2;152;130;179m \033[48;2;150;131;180m \033[48;2;148;132;181m \033[48;2;146;133;181m \033[48;2;140;130;177m \033[48;2;51;53;78m \033[48;2;54;57;81m \033[48;2;61;65;90m \033[48;2;54;60;84m \033[48;2;38;44;70m \033[48;2;44;51;77m \033[48;2;130;142;188m \033[48;2;128;143;189m \033[48;2;126;144;189m \033[48;2;125;146;191m \033[48;2;189;191;232m \033[48;2;120;147;192m \033[48;2;118;148;192m \033[48;2;116;149;193m \033[48;2;115;150;194m \033[48;2;113;150;194m \033[48;2;221;227;253m \033[48;2;223;227;252m \033[48;2;231;228;253m \033[48;2;237;223;248m \033[48;2;152;107;130m \033[48;2;184;102;131m \033[48;2;103;156;198m \033[48;2;103;156;199m \033[48;2;102;157;199m \033[48;2;101;157;199m \033[48;2;100;157;200m \033[48;2;106;83;129m \033[48;2;53;34;73m \033[48;2;203;199;236m \033[48;2;189;188;230m \033[48;2;187;187;223m \033[48;2;218;220;236m \033[48;2;255;255;255m \033[48;2;253;253;253m \033[48;2;254;254;254m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;118;151;194m \033[48;2;118;148;192m \033[48;2;120;147;192m \033[48;2;122;146;191m \033[48;2;124;145;190m \033[48;2;125;143;185m \033[48;2;21;24;31m \033[48;2;20;20;28m \033[48;2;21;18;27m \033[48;2;17;14;23m \033[48;2;16;11;18m \033[48;2;25;20;27m \033[48;2;32;27;34m \033[48;2;44;39;46m \033[48;2;44;40;46m \033[48;2;42;39;46m \033[48;2;44;39;46m \033[48;2;43;38;45m \033[48;2;41;34;42m \033[48;2;39;31;41m \033[48;2;39;31;42m \033[48;2;38;33;40m \033[48;2;37;32;39m \033[48;2;36;31;37m \033[48;2;34;29;33m \033[48;2;165;123;173m \033[48;2;167;122;173m \033[48;2;168;121;172m \033[48;2;170;120;171m \033[48;2;28;20;18m \033[48;2;32;21;19m \033[48;2;65;54;52m \033[48;2;80;65;65m \033[48;2;91;72;74m \033[48;2;62;46;49m \033[48;2;60;43;49m \033[48;2;46;32;39m \033[48;2;28;19;22m \033[48;2;20;12;11m \033[48;2;12;7;3m \033[48;2;13;8;4m \033[48;2;13;9;8m \033[m");
$display("\033[48;2;42;41;46m \033[48;2;44;43;49m \033[48;2;43;42;47m \033[48;2;45;44;50m \033[48;2;44;45;52m \033[48;2;47;47;55m \033[48;2;44;47;54m \033[48;2;44;47;54m \033[48;2;44;47;54m \033[48;2;44;47;54m \033[48;2;43;47;53m \033[48;2;172;120;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;167;122;173m \033[48;2;50;51;63m \033[48;2;45;49;58m \033[48;2;50;54;62m \033[48;2;50;54;63m \033[48;2;51;55;66m \033[48;2;51;54;69m \033[48;2;51;54;71m \033[48;2;151;130;179m \033[48;2;149;131;180m \033[48;2;147;132;181m \033[48;2;145;133;181m \033[48;2;48;52;77m \033[48;2;50;55;81m \033[48;2;53;58;84m \033[48;2;63;66;97m \033[48;2;56;59;90m \033[48;2;35;38;70m \033[48;2;131;141;187m \033[48;2;129;142;188m \033[48;2;127;143;189m \033[48;2;125;144;190m \033[48;2;206;207;251m \033[48;2;189;192;233m \033[48;2;197;199;240m \033[48;2;118;148;193m \033[48;2;116;149;193m \033[48;2;114;150;194m \033[48;2;112;151;195m \033[48;2;222;223;251m \033[48;2;226;226;249m \033[48;2;97;88;114m \033[48;2;106;80;108m \033[48;2;150;89;117m \033[48;2;186;98;120m \033[48;2;203;101;123m \033[48;2;101;157;199m \033[48;2;100;157;200m \033[48;2;99;158;200m \033[48;2;99;158;200m \033[48;2;98;158;201m \033[48;2;98;158;200m \033[48;2;99;158;200m \033[48;2;100;157;200m \033[48;2;103;158;200m \033[48;2;248;249;254m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;254;254;254m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;117;148;193m \033[48;2;119;147;192m \033[48;2;121;146;191m \033[48;2;123;145;190m \033[48;2;125;144;190m \033[48;2;127;143;189m \033[48;2;129;142;188m \033[48;2;131;141;187m \033[48;2;133;140;186m \033[48;2;32;22;29m \033[48;2;38;28;37m \033[48;2;46;37;48m \033[48;2;52;46;53m \033[48;2;52;46;53m \033[48;2;49;43;53m \033[48;2;47;41;51m \033[48;2;46;38;49m \033[48;2;45;37;48m \033[48;2;45;37;48m \033[48;2;44;36;48m \033[48;2;43;36;44m \033[48;2;41;33;41m \033[48;2;38;31;37m \033[48;2;36;31;36m \033[48;2;165;123;174m \033[48;2;166;122;173m \033[48;2;168;121;172m \033[48;2;170;120;171m \033[48;2;27;19;17m \033[48;2;30;20;18m \033[48;2;50;40;37m \033[48;2;78;64;63m \033[48;2;72;50;52m \033[48;2;69;44;47m \033[48;2;65;45;46m \033[48;2;61;45;45m \033[48;2;46;35;32m \033[48;2;22;12;8m \033[48;2;12;3;0m \033[48;2;14;5;2m \033[48;2;16;7;4m \033[m");
$display("\033[48;2;47;46;51m \033[48;2;48;47;53m \033[48;2;48;49;53m \033[48;2;48;49;54m \033[48;2;47;50;56m \033[48;2;47;50;57m \033[48;2;48;51;58m \033[48;2;48;51;58m \033[48;2;46;49;56m \033[48;2;48;51;58m \033[48;2;50;53;60m \033[48;2;172;120;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;167;122;173m \033[48;2;54;54;65m \033[48;2;49;52;61m \033[48;2;53;56;65m \033[48;2;54;57;66m \033[48;2;55;58;67m \033[48;2;151;125;173m \033[48;2;153;129;178m \033[48;2;151;130;179m \033[48;2;149;131;180m \033[48;2;147;132;181m \033[48;2;145;133;181m \033[48;2;52;54;77m \033[48;2;54;57;82m \033[48;2;60;65;91m \033[48;2;65;68;98m \033[48;2;64;67;98m \033[48;2;123;130;174m \033[48;2;131;141;187m \033[48;2;129;142;188m \033[48;2;127;143;189m \033[48;2;99;109;154m \033[48;2;147;148;192m \033[48;2;206;208;249m \033[48;2;203;206;247m \033[48;2;132;157;201m \033[48;2;116;149;193m \033[48;2;114;150;194m \033[48;2;112;151;195m \033[48;2;111;152;195m \033[48;2;5;4;35m \033[48;2;52;25;51m \033[48;2;93;37;66m \033[48;2;119;67;94m \033[48;2;122;84;129m \033[48;2;125;102;162m \033[48;2;136;102;157m \033[48;2;159;99;134m \033[48;2;99;158;200m \033[48;2;98;158;201m \033[48;2;97;159;201m \033[48;2;98;158;201m \033[48;2;99;158;200m \033[48;2;100;157;200m \033[48;2;101;157;199m \033[48;2;102;156;199m \033[48;2;103;156;198m \033[48;2;105;155;198m \033[48;2;150;183;213m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;121;146;191m \033[48;2;123;145;190m \033[48;2;125;144;190m \033[48;2;127;143;189m \033[48;2;129;142;188m \033[48;2;131;141;187m \033[48;2;133;140;187m \033[48;2;135;139;186m \033[48;2;137;138;185m \033[48;2;139;137;184m \033[48;2;141;136;183m \033[48;2;52;50;55m \033[48;2;53;48;55m \033[48;2;51;46;53m \033[48;2;50;43;51m \033[48;2;46;39;47m \033[48;2;45;37;48m \033[48;2;45;37;48m \033[48;2;44;37;45m \033[48;2;43;36;44m \033[48;2;38;31;39m \033[48;2;34;29;33m \033[48;2;165;123;174m \033[48;2;166;122;173m \033[48;2;168;121;172m \033[48;2;170;120;171m \033[48;2;28;18;16m \033[48;2;30;19;17m \033[48;2;31;19;15m \033[48;2;82;67;64m \033[48;2;59;37;35m \033[48;2;71;45;46m \033[48;2;70;44;44m \033[48;2;70;46;45m \033[48;2;55;31;31m \033[48;2;47;24;23m \033[48;2;46;22;22m \033[48;2;51;31;29m \033[48;2;50;31;27m \033[m");
$display("\033[48;2;50;49;54m \033[48;2;50;49;55m \033[48;2;48;51;55m \033[48;2;49;52;57m \033[48;2;47;50;55m \033[48;2;48;51;56m \033[48;2;50;53;60m \033[48;2;50;53;60m \033[48;2;51;54;61m \033[48;2;53;56;63m \033[48;2;55;58;65m \033[48;2;172;119;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;167;122;173m \033[48;2;165;123;173m \033[48;2;163;124;174m \033[48;2;161;125;175m \033[48;2;159;126;176m \033[48;2;157;127;177m \033[48;2;155;128;177m \033[48;2;154;129;178m \033[48;2;151;130;179m \033[48;2;150;131;180m \033[48;2;53;54;72m \033[48;2;52;53;73m \033[48;2;51;52;75m \033[48;2;58;60;84m \033[48;2;66;67;94m \033[48;2;65;68;99m \033[48;2;65;68;99m \033[48;2;133;140;186m \033[48;2;131;141;187m \033[48;2;129;142;188m \033[48;2;127;143;189m \033[48;2;72;74;115m \033[48;2;74;75;118m \033[48;2;165;167;210m \033[48;2;203;205;246m \033[48;2;208;210;249m \033[48;2;116;149;193m \033[48;2;115;150;194m \033[48;2;113;151;195m \033[48;2;111;151;195m \033[48;2;84;91;130m \033[48;2;17;3;30m \033[48;2;60;21;45m \033[48;2;87;34;58m \033[48;2;108;65;106m \033[48;2;119;94;157m \033[48;2;127;99;157m \033[48;2;140;100;147m \033[48;2;159;101;126m \033[48;2;118;57;83m \033[48;2;195;166;172m \033[48;2;251;250;255m \033[48;2;196;215;233m \033[48;2;101;157;199m \033[48;2;102;156;199m \033[48;2;103;156;199m \033[48;2;104;155;198m \033[48;2;105;155;198m \033[48;2;107;154;197m \033[48;2;108;153;196m \033[48;2;253;255;253m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;254m \033[48;2;252;255;255m \033[48;2;252;255;255m \033[48;2;254;255;255m \033[48;2;254;254;255m \033[48;2;253;254;253m \033[48;2;252;253;249m \033[48;2;248;247;237m \033[48;2;131;141;187m \033[48;2;133;140;186m \033[48;2;135;139;186m \033[48;2;137;138;185m \033[48;2;139;137;184m \033[48;2;141;136;183m \033[48;2;143;135;182m \033[48;2;58;51;60m \033[48;2;52;45;52m \033[48;2;53;46;50m \033[48;2;48;42;46m \033[48;2;46;39;46m \033[48;2;45;38;45m \033[48;2;45;38;45m \033[48;2;47;41;45m \033[48;2;38;32;36m \033[48;2;25;14;18m \033[48;2;165;123;174m \033[48;2;167;122;173m \033[48;2;168;121;172m \033[48;2;170;120;171m \033[48;2;29;19;17m \033[48;2;30;16;13m \033[48;2;34;20;17m \033[48;2;80;62;55m \033[48;2;72;50;38m \033[48;2;81;53;40m \033[48;2;82;50;38m \033[48;2;76;44;31m \033[48;2;71;41;30m \033[48;2;68;38;27m \033[48;2;66;38;26m \033[48;2;67;39;28m \033[48;2;66;39;30m \033[m");
$display("\033[48;2;52;51;56m \033[48;2;50;51;55m \033[48;2;50;52;57m \033[48;2;52;54;59m \033[48;2;51;54;59m \033[48;2;52;55;60m \033[48;2;53;56;63m \033[48;2;53;56;63m \033[48;2;53;56;63m \033[48;2;55;58;65m \033[48;2;57;59;67m \033[48;2;172;119;171m \033[48;2;170;120;171m \033[48;2;169;121;172m \033[48;2;167;122;173m \033[48;2;165;123;173m \033[48;2;164;124;174m \033[48;2;162;125;175m \033[48;2;147;117;163m \033[48;2;92;84;106m \033[48;2;58;61;70m \033[48;2;58;60;72m \033[48;2;56;58;71m \033[48;2;55;57;70m \033[48;2;53;54;74m \033[48;2;52;53;74m \033[48;2;51;53;77m \033[48;2;58;59;88m \033[48;2;66;67;97m \033[48;2;67;70;103m \033[48;2;136;138;185m \033[48;2;134;139;186m \033[48;2;132;141;187m \033[48;2;130;142;188m \033[48;2;128;143;188m \033[48;2;126;144;189m \033[48;2;124;145;190m \033[48;2;122;146;191m \033[48;2;121;146;191m \033[48;2;119;147;192m \033[48;2;117;148;193m \033[48;2;115;149;194m \033[48;2;114;150;194m \033[48;2;112;151;195m \033[48;2;111;152;195m \033[48;2;103;95;134m \033[48;2;59;33;68m \033[48;2;135;94;121m \033[48;2;159;108;146m \033[48;2;156;103;150m \033[48;2;165;103;143m \033[48;2;162;107;141m \033[48;2;170;109;140m \033[48;2;120;73;102m \033[48;2;230;209;217m \033[48;2;151;139;133m \033[48;2;248;239;233m \033[48;2;254;255;253m \033[48;2;254;255;253m \033[48;2;255;255;251m \033[48;2;106;155;198m \033[48;2;107;154;197m \033[48;2;108;153;197m \033[48;2;109;153;196m \033[48;2;111;152;195m \033[48;2;255;255;255m \033[48;2;255;255;255m \033[48;2;255;255;253m \033[48;2;255;255;253m \033[48;2;255;255;253m \033[48;2;255;255;252m \033[48;2;255;254;250m \033[48;2;252;253;248m \033[48;2;251;250;245m \033[48;2;213;207;182m \033[48;2;208;203;146m \033[48;2;92;87;39m \033[48;2;50;45;40m \033[48;2;45;43;48m \033[48;2;138;137;184m \033[48;2;140;136;184m \033[48;2;142;135;183m \033[48;2;144;134;182m \033[48;2;146;133;181m \033[48;2;52;45;52m \033[48;2;52;45;50m \033[48;2;53;47;51m \033[48;2;52;46;49m \033[48;2;49;43;47m \033[48;2;48;42;46m \033[48;2;48;42;46m \033[48;2;33;26;31m \033[48;2;12;2;8m \033[48;2;162;120;169m \033[48;2;167;122;173m \033[48;2;169;121;172m \033[48;2;170;120;171m \033[48;2;28;18;17m \033[48;2;31;17;14m \033[48;2;32;17;13m \033[48;2;74;56;49m \033[48;2;98;72;60m \033[48;2;104;70;53m \033[48;2;100;63;45m \033[48;2;98;62;46m \033[48;2;96;64;47m \033[48;2;89;57;40m \033[48;2;79;46;31m \033[48;2;78;46;31m \033[48;2;77;46;33m \033[m");
$display("\033[48;2;55;54;59m \033[48;2;55;55;60m \033[48;2;53;56;61m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;53;56;61m \033[48;2;53;56;63m \033[48;2;55;58;65m \033[48;2;57;59;66m \033[48;2;59;62;69m \033[48;2;61;64;71m \033[48;2;173;119;170m \033[48;2;171;120;171m \033[48;2;169;121;172m \033[48;2;168;122;172m \033[48;2;59;59;69m \033[48;2;55;58;65m \033[48;2;56;59;66m \033[48;2;56;59;66m \033[48;2;57;60;67m \033[48;2;55;57;69m \033[48;2;54;56;68m \033[48;2;54;56;69m \033[48;2;53;55;68m \033[48;2;53;54;75m \033[48;2;52;52;76m \033[48;2;52;52;80m \033[48;2;59;60;91m \033[48;2;73;73;107m \033[48;2;74;76;114m \033[48;2;137;138;185m \033[48;2;135;139;186m \033[48;2;133;140;186m \033[48;2;131;141;187m \033[48;2;129;142;188m \033[48;2;127;143;189m \033[48;2;125;144;189m \033[48;2;124;145;190m \033[48;2;122;146;191m \033[48;2;120;147;192m \033[48;2;118;148;192m \033[48;2;117;149;193m \033[48;2;115;149;194m \033[48;2;114;150;194m \033[48;2;112;151;195m \033[48;2;111;152;195m \033[48;2;110;93;133m \033[48;2;127;91;140m \033[48;2;168;110;153m \033[48;2;181;106;133m \033[48;2;201;106;116m \033[48;2;200;108;120m \033[48;2;187;99;128m \033[48;2;123;76;105m \033[48;2;203;182;208m \033[48;2;114;90;64m \033[48;2;129;85;26m \033[48;2;157;121;62m \033[48;2;242;215;168m \033[48;2;208;188;144m \033[48;2;107;153;197m \033[48;2;109;153;196m \033[48;2;110;152;196m \033[48;2;111;152;195m \033[48;2;185;204;224m \033[48;2;255;255;253m \033[48;2;255;255;253m \033[48;2;255;255;250m \033[48;2;241;242;237m \033[48;2;212;208;197m \033[48;2;224;218;201m \033[48;2;189;177;151m \033[48;2;181;165;129m \033[48;2;233;214;172m \033[48;2;146;124;69m \033[48;2;132;109;47m \033[48;2;67;49;30m \033[48;2;50;46;58m \033[48;2;45;44;50m \033[48;2;139;137;184m \033[48;2;141;136;183m \033[48;2;143;135;182m \033[48;2;145;134;182m \033[48;2;147;133;181m \033[48;2;57;50;57m \033[48;2;54;48;53m \033[48;2;54;48;52m \033[48;2;54;48;52m \033[48;2;54;48;52m \033[48;2;51;45;49m \033[48;2;41;35;39m \033[48;2;11;5;9m \033[48;2;32;24;32m \033[48;2;46;40;44m \033[48;2;39;33;35m \033[48;2;25;19;21m \033[48;2;25;15;13m \033[48;2;27;17;16m \033[48;2;33;19;16m \033[48;2;32;18;15m \033[48;2;40;23;15m \033[48;2;102;73;58m \033[48;2;106;69;51m \033[48;2;101;61;41m \033[48;2;99;60;40m \033[48;2;94;54;34m \033[48;2;77;40;18m \033[48;2;79;41;22m \033[48;2;71;34;14m \033[48;2;74;38;21m \033[m");
$display("\033[48;2;55;55;57m \033[48;2;55;56;58m \033[48;2;53;56;61m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;55;58;65m \033[48;2;56;59;66m \033[48;2;58;61;68m \033[48;2;59;62;69m \033[48;2;61;64;69m \033[48;2;173;119;170m \033[48;2;171;120;171m \033[48;2;170;120;171m \033[48;2;168;121;172m \033[48;2;59;59;69m \033[48;2;55;58;67m \033[48;2;55;58;67m \033[48;2;56;58;70m \033[48;2;58;60;72m \033[48;2;55;57;72m \033[48;2;53;54;72m \033[48;2;53;54;74m \033[48;2;52;53;74m \033[48;2;55;53;77m \033[48;2;53;53;79m \033[48;2;54;53;84m \033[48;2;60;60;95m \033[48;2;73;73;112m \033[48;2;140;136;184m \033[48;2;138;137;184m \033[48;2;136;138;185m \033[48;2;134;139;186m \033[48;2;70;73;116m \033[48;2;71;74;119m \033[48;2;74;77;125m \033[48;2;71;75;124m \033[48;2;75;78;129m \033[48;2;76;78;127m \033[48;2;75;77;125m \033[48;2;185;190;231m \033[48;2;206;211;251m \033[48;2;117;148;193m \033[48;2;116;149;193m \033[48;2;114;150;194m \033[48;2;113;150;194m \033[48;2;123;117;165m \033[48;2;101;70;118m \033[48;2;162;105;150m \033[48;2;109;153;196m \033[48;2;108;153;196m \033[48;2;108;153;197m \033[48;2;107;154;197m \033[48;2;107;154;197m \033[48;2;107;154;197m \033[48;2;107;154;197m \033[48;2;107;154;197m \033[48;2;108;153;197m \033[48;2;108;153;196m \033[48;2;109;153;196m \033[48;2;110;152;196m \033[48;2;111;152;195m \033[48;2;112;151;195m \033[48;2;113;151;194m \033[48;2;211;201;158m \033[48;2;192;177;114m \033[48;2;244;232;181m \033[48;2;252;244;200m \033[48;2;120;147;192m \033[48;2;122;146;191m \033[48;2;123;145;190m \033[48;2;125;144;190m \033[48;2;127;143;189m \033[48;2;129;142;188m \033[48;2;131;141;187m \033[48;2;132;140;187m \033[48;2;134;139;186m \033[48;2;136;138;185m \033[48;2;138;137;184m \033[48;2;140;136;184m \033[48;2;142;135;183m \033[48;2;144;134;182m \033[48;2;146;133;181m \033[48;2;57;55;60m \033[48;2;55;50;56m \033[48;2;55;50;55m \033[48;2;56;50;54m \033[48;2;56;50;54m \033[48;2;55;49;53m \033[48;2;54;48;52m \033[48;2;31;25;29m \033[48;2;23;17;21m \033[48;2;46;39;44m \033[48;2;166;122;173m \033[48;2;168;121;172m \033[48;2;170;121;172m \033[48;2;171;120;171m \033[48;2;173;119;170m \033[48;2;17;9;7m \033[48;2;17;10;4m \033[48;2;19;9;3m \033[48;2;12;1;1m \033[48;2;28;8;3m \033[48;2;71;46;36m \033[48;2;124;92;82m \033[48;2;148;112;94m \033[48;2;138;101;81m \033[48;2;136;94;72m \033[48;2;132;88;64m \033[48;2;127;82;57m \033[m");
$display("\033[48;2;56;56;58m \033[48;2;56;57;59m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;53;56;61m \033[48;2;54;57;63m \033[48;2;59;62;67m \033[48;2;58;61;65m \033[48;2;60;63;68m \033[48;2;62;65;70m \033[48;2;174;118;170m \033[48;2;172;119;171m \033[48;2;171;120;171m \033[48;2;169;121;172m \033[48;2;58;58;69m \033[48;2;53;55;67m \033[48;2;54;56;69m \033[48;2;55;57;70m \033[48;2;56;58;71m \033[48;2;54;56;69m \033[48;2;53;55;70m \033[48;2;52;53;71m \033[48;2;52;53;73m \033[48;2;53;53;79m \033[48;2;52;53;81m \033[48;2;53;53;87m \033[48;2;58;61;97m \033[48;2;117;113;157m \033[48;2;141;136;183m \033[48;2;139;136;184m \033[48;2;138;137;185m \033[48;2;136;138;185m \033[48;2;65;63;103m \033[48;2;68;70;111m \033[48;2;74;74;118m \033[48;2;73;76;121m \033[48;2;73;76;121m \033[48;2;74;77;120m \033[48;2;77;80;123m \033[48;2;77;82;124m \033[48;2;121;126;166m \033[48;2;119;147;192m \033[48;2;118;148;192m \033[48;2;117;149;193m \033[48;2;116;149;193m \033[48;2;115;150;194m \033[48;2;94;47;76m \033[48;2;181;110;139m \033[48;2;112;151;195m \033[48;2;111;151;195m \033[48;2;111;152;195m \033[48;2;110;152;196m \033[48;2;110;152;196m \033[48;2;110;152;196m \033[48;2;110;152;196m \033[48;2;110;152;196m \033[48;2;111;152;195m \033[48;2;111;151;195m \033[48;2;112;151;195m \033[48;2;113;151;195m \033[48;2;114;150;194m \033[48;2;245;213;127m \033[48;2;238;215;134m \033[48;2;192;176;107m \033[48;2;207;199;128m \033[48;2;242;239;186m \033[48;2;246;248;203m \033[48;2;122;146;191m \033[48;2;124;145;190m \033[48;2;125;144;190m \033[48;2;127;143;189m \033[48;2;129;142;188m \033[48;2;130;141;187m \033[48;2;132;140;187m \033[48;2;134;139;186m \033[48;2;136;138;185m \033[48;2;138;138;185m \033[48;2;139;137;184m \033[48;2;141;136;183m \033[48;2;143;135;182m \033[48;2;54;51;58m \033[48;2;57;54;61m \033[48;2;56;54;57m \033[48;2;57;52;56m \033[48;2;56;52;53m \033[48;2;58;52;54m \033[48;2;57;51;53m \033[48;2;59;53;55m \033[48;2;51;45;47m \033[48;2;30;24;26m \033[48;2;49;43;46m \033[48;2;33;26;33m \033[48;2;167;122;173m \033[48;2;169;121;172m \033[48;2;171;120;171m \033[48;2;172;119;171m \033[48;2;159;108;155m \033[48;2;6;1;5m \033[48;2;5;1;5m \033[48;2;3;1;6m \033[48;2;2;2;7m \033[48;2;4;5;9m \033[48;2;14;9;15m \033[48;2;16;12;20m \033[48;2;13;11;18m \033[48;2;18;11;21m \033[48;2;23;12;22m \033[48;2;20;7;16m \033[48;2;22;6;13m \033[m");
$display("\033[48;2;58;58;60m \033[48;2;57;58;59m \033[48;2;55;58;63m \033[48;2;55;58;63m \033[48;2;55;58;63m \033[48;2;55;58;63m \033[48;2;59;62;67m \033[48;2;60;63;68m \033[48;2;61;64;69m \033[48;2;61;64;69m \033[48;2;62;65;70m \033[48;2;63;66;71m \033[48;2;65;68;73m \033[48;2;42;45;50m \033[48;2;46;49;54m \033[48;2;48;50;59m \033[48;2;53;56;65m \033[48;2;53;57;68m \033[48;2;53;57;68m \033[48;2;53;57;68m \033[48;2;53;57;68m \033[48;2;53;57;68m \033[48;2;51;54;69m \033[48;2;51;54;73m \033[48;2;51;53;74m \033[48;2;52;54;77m \033[48;2;49;53;82m \033[48;2;62;65;97m \033[48;2;77;81;116m \033[48;2;72;74;112m \033[48;2;57;59;97m \033[48;2;55;57;95m \033[48;2;56;58;96m \033[48;2;60;63;104m \033[48;2;61;63;105m \033[48;2;60;64;103m \033[48;2;63;67;105m \033[48;2;70;74;112m \033[48;2;74;78;116m \033[48;2;76;79;119m \033[48;2;75;80;121m \033[48;2;80;85;126m \033[48;2;117;125;169m \033[48;2;132;144;185m \033[48;2;99;100;134m \033[48;2;119;67;96m \033[48;2;183;90;116m \033[48;2;115;29;51m \033[48;2;200;106;131m \033[48;2;178;96;131m \033[48;2;133;96;151m \033[48;2;101;88;153m \033[48;2;114;81;140m \033[48;2;115;70;109m \033[48;2;103;54;86m \033[48;2;134;88;64m \033[48;2;156;109;41m \033[48;2;202;157;63m \033[48;2;225;185;89m \033[48;2;224;188;92m \033[48;2;205;175;71m \033[48;2;224;194;98m \033[48;2;223;202;123m \033[48;2;249;240;179m \033[48;2;255;244;192m \033[48;2;254;244;185m \033[48;2;233;225;167m \033[48;2;231;222;164m \033[48;2;241;226;168m \033[48;2;239;222;160m \033[48;2;239;221;153m \033[48;2;250;230;156m \033[48;2;177;154;79m \033[48;2;198;173;98m \033[48;2;121;91;45m \033[48;2;72;55;51m \033[48;2;59;56;67m \033[48;2;62;58;64m \033[48;2;56;55;63m \033[48;2;57;54;63m \033[48;2;56;53;60m \033[48;2;59;54;61m \033[48;2;60;55;61m \033[48;2;59;54;60m \033[48;2;57;52;56m \033[48;2;55;50;54m \033[48;2;57;53;56m \033[48;2;60;54;56m \033[48;2;59;53;55m \033[48;2;37;31;33m \033[48;2;38;32;34m \033[48;2;34;28;30m \033[48;2;14;8;10m \033[48;2;19;13;15m \033[48;2;30;24;28m \033[48;2;29;23;27m \033[48;2;32;27;31m \033[48;2;4;0;3m \033[48;2;2;0;3m \033[48;2;2;0;3m \033[48;2;1;1;3m \033[48;2;1;0;4m \033[48;2;1;0;4m \033[48;2;1;0;6m \033[48;2;2;1;6m \033[48;2;2;2;8m \033[48;2;2;2;10m \033[48;2;0;1;10m \033[48;2;0;2;12m \033[48;2;2;4;13m \033[m");
$display("\033[48;2;59;59;61m \033[48;2;57;58;60m \033[48;2;56;59;64m \033[48;2;56;58;63m \033[48;2;55;58;63m \033[48;2;58;61;66m \033[48;2;61;63;68m \033[48;2;61;64;69m \033[48;2;63;66;72m \033[48;2;65;68;73m \033[48;2;66;68;74m \033[48;2;65;68;73m \033[48;2;66;69;74m \033[48;2;55;58;63m \033[48;2;54;57;62m \033[48;2;46;49;56m \033[48;2;51;55;61m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;52;56;67m \033[48;2;51;54;69m \033[48;2;52;54;75m \033[48;2;54;56;79m \033[48;2;53;57;86m \033[48;2;62;65;97m \033[48;2;73;77;113m \033[48;2;71;73;112m \033[48;2;51;53;92m \033[48;2;63;65;104m \033[48;2;59;61;100m \033[48;2;61;63;105m \033[48;2;60;63;104m \033[48;2;60;64;102m \033[48;2;60;64;102m \033[48;2;66;69;107m \033[48;2;69;73;110m \033[48;2;71;75;112m \033[48;2;73;79;113m \033[48;2;77;83;115m \033[48;2;90;96;130m \033[48;2;145;149;187m \033[48;2;54;51;82m \033[48;2;122;74;98m \033[48;2;169;83;106m \033[48;2;95;23;57m \033[48;2;154;92;128m \033[48;2;155;89;111m \033[48;2;157;84;100m \033[48;2;157;77;95m \033[48;2;148;73;89m \033[48;2;129;78;112m \033[48;2;107;73;114m \033[48;2;108;73;48m \033[48;2;157;107;41m \033[48;2;182;133;44m \033[48;2;200;154;62m \033[48;2;198;157;64m \033[48;2;242;205;108m \033[48;2;249;218;130m \033[48;2;248;221;146m \033[48;2;239;217;150m \033[48;2;248;231;165m \033[48;2;236;215;148m \033[48;2;220;200;133m \033[48;2;229;211;144m \033[48;2;246;232;162m \033[48;2;239;218;153m \033[48;2;244;219;149m \033[48;2;243;211;135m \033[48;2;251;216;136m \033[48;2;223;187;112m \033[48;2;94;72;29m \033[48;2;75;64;64m \033[48;2;67;64;72m \033[48;2;66;63;71m \033[48;2;58;57;65m \033[48;2;56;53;62m \033[48;2;59;56;63m \033[48;2;64;59;65m \033[48;2;61;56;62m \033[48;2;58;53;59m \033[48;2;54;49;53m \033[48;2;57;52;56m \033[48;2;60;56;59m \033[48;2;62;56;58m \033[48;2;54;48;50m \033[48;2;37;31;33m \033[48;2;27;21;23m \033[48;2;21;15;17m \033[48;2;42;36;38m \033[48;2;40;34;36m \033[48;2;35;29;33m \033[48;2;34;28;32m \033[48;2;37;32;36m \033[48;2;2;0;1m \033[48;2;2;0;3m \033[48;2;2;0;3m \033[48;2;1;1;3m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[48;2;1;0;2m \033[48;2;0;0;4m \033[48;2;1;0;5m \033[48;2;0;1;6m \033[48;2;0;1;6m \033[m");
$display("\033[48;2;61;60;66m \033[48;2;62;60;66m \033[48;2;60;61;66m \033[48;2;57;60;65m \033[48;2;57;60;65m \033[48;2;62;66;71m \033[48;2;63;68;72m \033[48;2;64;69;73m \033[48;2;64;69;73m \033[48;2;64;69;73m \033[48;2;64;69;73m \033[48;2;65;70;74m \033[48;2;65;70;74m \033[48;2;59;64;68m \033[48;2;39;44;48m \033[48;2;48;52;62m \033[48;2;52;56;65m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;53;57;66m \033[48;2;55;57;69m \033[48;2;55;57;69m \033[48;2;54;56;69m \033[48;2;53;55;68m \033[48;2;54;57;74m \033[48;2;57;59;80m \033[48;2;57;62;89m \033[48;2;65;70;104m \033[48;2;75;79;119m \033[48;2;77;84;125m \033[48;2;52;56;101m \033[48;2;67;71;117m \033[48;2;72;75;123m \033[48;2;69;74;122m \033[48;2;68;70;117m \033[48;2;62;65;107m \033[48;2;60;63;100m \033[48;2;63;66;101m \033[48;2;67;70;103m \033[48;2;70;73;104m \033[48;2;72;76;105m \033[48;2;75;78;107m \033[48;2;75;80;109m \033[48;2;72;75;102m \033[48;2;57;51;79m \033[48;2;82;61;92m \033[48;2;88;58;89m \033[48;2;50;15;49m \033[48;2;123;89;131m \033[48;2;142;87;114m \033[48;2;164;77;89m \033[48;2;152;64;82m \033[48;2;158;67;80m \033[48;2;133;75;111m \033[48;2;119;87;118m \033[48;2;133;93;79m \033[48;2;140;87;23m \033[48;2;187;136;55m \033[48;2;239;199;123m \033[48;2;250;223;149m \033[48;2;236;208;127m \033[48;2;230;198;116m \033[48;2;233;204;124m \033[48;2;242;221;147m \033[48;2;252;237;167m \033[48;2;244;235;164m \033[48;2;255;245;178m \033[48;2;253;232;165m \033[48;2;243;214;145m \033[48;2;237;205;131m \033[48;2;238;203;124m \033[48;2;227;179;103m \033[48;2;211;164;80m \033[48;2;153;118;60m \033[48;2;81;68;52m \033[48;2;69;66;81m \033[48;2;69;65;77m \033[48;2;62;61;70m \033[48;2;60;58;69m \033[48;2;55;53;64m \033[48;2;61;59;70m \033[48;2;62;60;71m \033[48;2;62;60;70m \033[48;2;59;55;65m \033[48;2;57;54;61m \033[48;2;60;55;61m \033[48;2;61;56;60m \033[48;2;62;56;58m \033[48;2;48;43;44m \033[48;2;25;19;21m \033[48;2;41;35;37m \033[48;2;45;39;41m \033[48;2;49;39;42m \033[48;2;43;34;37m \033[48;2;35;29;33m \033[48;2;24;18;22m \033[48;2;15;11;15m \033[48;2;6;4;7m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;1;1;2m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[48;2;0;0;2m \033[m");
$display("\033[48;2;61;60;66m \033[48;2;60;61;66m \033[48;2;58;61;66m \033[48;2;57;62;66m \033[48;2;59;64;68m \033[48;2;64;69;73m \033[48;2;62;70;73m \033[48;2;63;71;74m \033[48;2;63;71;74m \033[48;2;64;72;75m \033[48;2;64;72;75m \033[48;2;64;72;75m \033[48;2;64;72;75m \033[48;2;66;74;77m \033[48;2;39;47;50m \033[48;2;48;52;61m \033[48;2;51;55;64m \033[48;2;52;56;65m \033[48;2;53;57;66m \033[48;2;54;58;67m \033[48;2;56;59;68m \033[48;2;57;59;71m \033[48;2;57;59;72m \033[48;2;58;60;73m \033[48;2;58;61;78m \033[48;2;59;61;82m \033[48;2;58;63;91m \033[48;2;65;70;104m \033[48;2;73;78;119m \033[48;2;75;82;126m \033[48;2;54;58;105m \033[48;2;66;70;117m \033[48;2;72;76;124m \033[48;2;72;75;128m \033[48;2;72;75;125m \033[48;2;72;75;120m \033[48;2;65;68;109m \033[48;2;66;68;106m \033[48;2;65;67;105m \033[48;2;66;69;102m \033[48;2;67;70;100m \033[48;2;68;72;98m \033[48;2;67;72;97m \033[48;2;70;74;101m \033[48;2;67;66;95m \033[48;2;41;31;65m \033[48;2;45;28;62m \033[48;2;33;9;45m \033[48;2;107;79;116m \033[48;2;108;65;96m \033[48;2;120;60;80m \033[48;2;123;57;77m \033[48;2;122;54;71m \033[48;2;119;56;77m \033[48;2;140;83;84m \033[48;2;143;87;57m \033[48;2;153;97;35m \033[48;2;217;159;75m \033[48;2;206;152;63m \033[48;2;230;185;94m \033[48;2;218;178;88m \033[48;2;202;166;80m \033[48;2;238;211;129m \033[48;2;252;233;154m \033[48;2;252;233;157m \033[48;2;240;214;142m \033[48;2;250;226;155m \033[48;2;235;207;136m \033[48;2;244;211;139m \033[48;2;244;210;139m \033[48;2;230;194;112m \033[48;2;224;177;97m \033[48;2;174;128;46m \033[48;2;103;71;20m \033[48;2;80;66;56m \033[48;2;68;65;80m \033[48;2;67;64;74m \033[48;2;58;57;68m \033[48;2;59;57;68m \033[48;2;58;56;67m \033[48;2;62;60;71m \033[48;2;64;62;73m \033[48;2;66;64;75m \033[48;2;63;62;69m \033[48;2;56;53;60m \033[48;2;62;57;63m \033[48;2;64;59;63m \033[48;2;61;55;57m \033[48;2;39;33;34m \033[48;2;18;12;14m \033[48;2;11;5;7m \033[48;2;9;2;4m \033[48;2;8;0;2m \033[48;2;8;0;2m \033[48;2;13;5;10m \033[48;2;27;20;25m \033[48;2;39;37;40m \033[48;2;28;26;29m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;1;1;2m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;0;0;0m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[48;2;1;1;3m \033[m");
$display ("----------------------------------------------------------------------------------------------------");
$display ("                                    Xian Zai Wo You Bing Qi Lin!                                    ");
$display ("----------------------------------------------------------------------------------------------------");
end endtask

task RickRoll; begin
$display("\033[48;2;168;153;186m \033[48;2;168;153;186m \033[48;2;168;153;186m \033[48;2;168;153;186m \033[48;2;168;153;186m \033[48;2;164;150;182m \033[48;2;165;152;180m \033[48;2;165;152;178m \033[48;2;165;152;178m \033[48;2;165;152;178m \033[48;2;161;148;174m \033[48;2;160;145;176m \033[48;2;160;145;176m \033[48;2;160;145;176m \033[48;2;162;148;174m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[48;2;163;147;174m \033[48;2;163;147;174m \033[48;2;163;147;174m \033[48;2;162;146;173m \033[48;2;161;145;171m \033[48;2;163;147;173m \033[48;2;163;147;173m \033[48;2;167;147;174m \033[48;2;166;146;173m \033[48;2;164;144;171m \033[48;2;164;144;171m \033[48;2;164;144;171m \033[48;2;164;144;171m \033[48;2;163;143;170m \033[48;2;166;146;171m \033[48;2;164;145;165m \033[48;2;163;143;166m \033[48;2;165;143;166m \033[48;2;167;141;166m \033[48;2;170;142;164m \033[48;2;170;142;159m \033[48;2;177;141;147m \033[48;2;183;132;128m \033[48;2;177;119;106m \033[48;2;167;104;76m \033[48;2;143;71;47m \033[48;2;116;51;27m \033[48;2;115;54;32m \033[48;2;108;58;33m \033[48;2;100;50;25m \033[48;2;93;44;22m \033[48;2;96;47;29m \033[48;2;97;51;31m \033[48;2;99;58;35m \033[48;2;97;51;36m \033[48;2;94;50;31m \033[48;2;91;47;23m \033[48;2;91;52;23m \033[48;2;96;57;34m \033[48;2;107;70;52m \033[48;2;113;75;62m \033[48;2;111;71;60m \033[48;2;110;67;55m \033[48;2;116;69;56m \033[48;2;112;65;53m \033[48;2;117;69;56m \033[48;2;122;74;64m \033[48;2;121;75;68m \033[48;2;121;76;77m \033[48;2;133;99;107m \033[48;2;173;143;158m \033[48;2;173;152;174m \033[48;2;170;150;177m \033[48;2;170;150;176m \033[48;2;173;153;179m \033[48;2;173;153;178m \033[48;2;173;153;178m \033[48;2;172;152;177m \033[48;2;173;153;178m \033[48;2;173;153;178m \033[48;2;170;150;175m \033[48;2;169;151;175m \033[48;2;167;151;175m \033[48;2;167;151;175m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;173m \033[48;2;166;152;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;163;149;174m \033[48;2;163;149;174m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;161;151;176m \033[48;2;162;153;174m \033[m");
$display("\033[48;2;171;158;189m \033[48;2;171;158;187m \033[48;2;171;158;189m \033[48;2;171;157;188m \033[48;2;171;157;188m \033[48;2;170;156;187m \033[48;2;169;156;186m \033[48;2;169;156;185m \033[48;2;169;156;182m \033[48;2;169;156;182m \033[48;2;167;154;180m \033[48;2;165;151;179m \033[48;2;165;151;178m \033[48;2;166;152;179m \033[48;2;169;155;181m \033[48;2;167;153;179m \033[48;2;167;153;179m \033[48;2;166;150;177m \033[48;2;166;150;177m \033[48;2;166;150;177m \033[48;2;165;149;176m \033[48;2;163;147;174m \033[48;2;163;147;174m \033[48;2;163;147;173m \033[48;2;163;147;173m \033[48;2;162;146;172m \033[48;2;164;146;172m \033[48;2;163;147;173m \033[48;2;164;147;173m \033[48;2;167;147;172m \033[48;2;167;147;172m \033[48;2;167;147;172m \033[48;2;166;148;173m \033[48;2;167;148;170m \033[48;2;168;146;166m \033[48;2;166;145;162m \033[48;2;173;145;154m \033[48;2;182;142;143m \033[48;2;184;140;135m \033[48;2;190;144;138m \033[48;2;192;140;131m \033[48;2;186;119;103m \033[48;2;159;90;68m \033[48;2;151;78;48m \033[48;2;141;69;38m \033[48;2;122;56;25m \033[48;2;118;55;31m \033[48;2;95;44;17m \033[48;2;88;42;16m \033[48;2;85;49;22m \033[48;2;83;47;27m \033[48;2;87;53;33m \033[48;2;91;56;39m \033[48;2;96;61;49m \033[48;2;98;65;51m \033[48;2;87;52;40m \033[48;2;94;58;44m \033[48;2;93;55;45m \033[48;2;102;62;56m \033[48;2;108;71;63m \033[48;2;99;61;54m \033[48;2;96;58;49m \033[48;2;92;56;40m \033[48;2;90;54;38m \033[48;2;102;66;50m \033[48;2;106;66;54m \033[48;2;110;71;63m \033[48;2;118;78;74m \033[48;2;123;84;84m \033[48;2;154;114;117m \033[48;2;181;143;159m \033[48;2;182;157;172m \033[48;2;175;157;173m \033[48;2;174;156;176m \033[48;2;175;155;180m \033[48;2;175;155;180m \033[48;2;174;154;179m \033[48;2;176;156;182m \033[48;2;176;156;182m \033[48;2;175;155;181m \033[48;2;173;154;183m \033[48;2;171;155;183m \033[48;2;170;154;181m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;166;152;178m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[48;2;164;149;180m \033[48;2;163;148;179m \033[48;2;164;149;180m \033[48;2;170;155;186m \033[48;2;171;155;183m \033[48;2;170;154;181m \033[48;2;165;149;177m \033[48;2;163;148;174m \033[48;2;164;149;175m \033[48;2;164;148;175m \033[48;2;163;149;174m \033[48;2;163;149;174m \033[48;2;164;150;176m \033[48;2;164;149;178m \033[48;2;164;149;178m \033[48;2;165;150;181m \033[48;2;164;151;180m \033[48;2;162;151;180m \033[48;2;163;153;180m \033[m");
$display("\033[48;2;176;163;193m \033[48;2;173;160;188m \033[48;2;172;159;189m \033[48;2;171;158;188m \033[48;2;170;157;187m \033[48;2;172;159;188m \033[48;2;172;159;189m \033[48;2;172;159;189m \033[48;2;169;156;182m \033[48;2;170;157;183m \033[48;2;166;153;179m \033[48;2;166;152;178m \033[48;2;167;153;179m \033[48;2;168;154;180m \033[48;2;169;155;181m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;167;151;178m \033[48;2;167;151;178m \033[48;2;167;151;178m \033[48;2;166;150;177m \033[48;2;164;148;175m \033[48;2;165;149;176m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;167;147;172m \033[48;2;167;147;172m \033[48;2;167;147;172m \033[48;2;168;148;168m \033[48;2;169;146;165m \033[48;2;171;146;161m \033[48;2;175;139;141m \033[48;2;184;140;130m \033[48;2;185;130;108m \033[48;2;177;111;81m \033[48;2;183;117;85m \033[48;2;173;103;68m \033[48;2;161;96;64m \033[48;2;157;89;57m \033[48;2;155;80;51m \033[48;2;137;72;37m \033[48;2;126;65;32m \033[48;2;115;59;34m \033[48;2;108;63;39m \033[48;2;87;50;26m \033[48;2;83;55;34m \033[48;2;83;54;30m \033[48;2;80;51;31m \033[48;2;86;56;38m \033[48;2;88;55;36m \033[48;2;85;53;33m \033[48;2;77;44;25m \033[48;2;87;52;33m \033[48;2;90;53;38m \033[48;2;94;58;46m \033[48;2;101;65;53m \033[48;2;96;60;45m \033[48;2;93;58;38m \033[48;2;91;55;39m \033[48;2;89;53;37m \033[48;2;90;54;38m \033[48;2;96;58;47m \033[48;2;98;59;51m \033[48;2;112;73;68m \033[48;2;113;74;68m \033[48;2;110;71;64m \033[48;2;118;77;76m \033[48;2;167;138;139m \033[48;2;178;157;164m \033[48;2;176;152;175m \033[48;2;177;155;180m \033[48;2;175;155;180m \033[48;2;175;155;180m \033[48;2;175;155;182m \033[48;2;175;155;182m \033[48;2;174;154;181m \033[48;2;174;156;183m \033[48;2;172;156;183m \033[48;2;171;155;182m \033[48;2;169;155;181m \033[48;2;169;155;181m \033[48;2;171;157;183m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;168;154;180m \033[48;2;165;151;180m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[48;2;168;153;184m \033[48;2;172;156;185m \033[48;2;172;156;183m \033[48;2;175;159;186m \033[48;2;170;154;181m \033[48;2;166;150;177m \033[48;2;165;149;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;149;179m \033[48;2;164;149;180m \033[48;2;165;150;181m \033[48;2;164;151;181m \033[48;2;162;151;181m \033[48;2;163;152;182m \033[m");
$display("\033[48;2;185;171;204m \033[48;2;182;168;201m \033[48;2;177;164;194m \033[48;2;186;173;203m \033[48;2;186;173;203m \033[48;2;183;173;198m \033[48;2;182;172;197m \033[48;2;179;169;194m \033[48;2;175;165;190m \033[48;2;176;166;191m \033[48;2;173;163;188m \033[48;2;170;162;185m \033[48;2;177;167;191m \033[48;2;180;166;189m \033[48;2;180;166;191m \033[48;2;176;162;187m \033[48;2;172;158;183m \033[48;2;171;157;183m \033[48;2;168;154;180m \033[48;2;168;154;180m \033[48;2;169;153;180m \033[48;2;167;151;177m \033[48;2;166;151;174m \033[48;2;165;150;173m \033[48;2;165;150;173m \033[48;2;165;150;173m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;149;172m \033[48;2;164;149;172m \033[48;2;164;149;172m \033[48;2;164;146;165m \033[48;2;170;144;157m \033[48;2;145;100;99m \033[48;2;163;110;91m \033[48;2;177;124;90m \033[48;2;172;116;76m \033[48;2;164;105;68m \033[48;2;165;105;69m \033[48;2;157;92;62m \033[48;2;153;84;52m \033[48;2;159;92;61m \033[48;2;147;82;50m \033[48;2;134;67;39m \033[48;2;120;63;38m \033[48;2;103;54;32m \033[48;2;89;51;30m \033[48;2;83;48;28m \033[48;2;88;55;38m \033[48;2;91;59;41m \033[48;2;88;56;37m \033[48;2;85;54;36m \033[48;2;80;50;28m \033[48;2;75;44;23m \033[48;2;78;46;25m \033[48;2;81;49;28m \033[48;2;86;54;33m \033[48;2;90;58;37m \033[48;2;92;58;38m \033[48;2;93;57;41m \033[48;2;94;58;45m \033[48;2;91;55;37m \033[48;2;95;59;42m \033[48;2;99;63;47m \033[48;2;95;57;45m \033[48;2;96;57;49m \033[48;2;112;73;68m \033[48;2;110;76;67m \033[48;2;124;81;75m \033[48;2;128;88;81m \033[48;2;154;122;118m \033[48;2;176;149;156m \033[48;2;176;153;170m \033[48;2;174;155;175m \033[48;2;174;155;177m \033[48;2;173;153;180m \033[48;2;169;153;179m \033[48;2;169;153;179m \033[48;2;167;151;177m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;169;155;181m \033[48;2;169;155;181m \033[48;2;169;155;181m \033[48;2;172;158;184m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;167;153;179m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;164;150;179m \033[48;2;165;150;181m \033[48;2;172;157;188m \033[48;2;172;156;187m \033[48;2;173;159;185m \033[48;2;169;155;181m \033[48;2;167;151;178m \033[48;2;167;151;178m \033[48;2;165;149;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;161;151;176m \033[48;2;163;151;179m \033[48;2;164;151;181m \033[48;2;164;151;181m \033[48;2;164;151;181m \033[48;2;163;152;182m \033[48;2;164;153;183m \033[m");
$display("\033[48;2;188;177;209m \033[48;2;186;175;207m \033[48;2;185;172;202m \033[48;2;182;169;199m \033[48;2;185;172;202m \033[48;2;185;172;202m \033[48;2;185;172;202m \033[48;2;186;172;203m \033[48;2;186;172;202m \033[48;2;185;171;202m \033[48;2;172;159;189m \033[48;2;172;159;185m \033[48;2;179;166;192m \033[48;2;179;167;192m \033[48;2;180;166;191m \033[48;2;184;170;195m \033[48;2;178;164;189m \033[48;2;172;158;184m \033[48;2;170;156;182m \033[48;2;169;155;181m \033[48;2;169;153;180m \033[48;2;167;151;178m \033[48;2;167;151;178m \033[48;2;166;151;173m \033[48;2;166;151;173m \033[48;2;166;151;173m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;148;174m \033[48;2;164;149;172m \033[48;2;164;149;170m \033[48;2;165;151;168m \033[48;2;172;153;164m \033[48;2;160;128;124m \033[48;2;176;134;111m \033[48;2;181;133;93m \033[48;2;191;135;96m \033[48;2;175;125;79m \033[48;2;169;115;84m \033[48;2;162;105;77m \033[48;2;148;89;64m \033[48;2;140;81;48m \033[48;2;137;76;48m \033[48;2;142;85;64m \033[48;2;130;82;58m \033[48;2;125;80;57m \033[48;2;122;77;58m \033[48;2;110;78;57m \033[48;2;111;76;63m \033[48;2;110;75;68m \033[48;2;109;69;65m \033[48;2;106;66;61m \033[48;2;98;59;54m \033[48;2;96;59;44m \033[48;2;96;59;44m \033[48;2;98;62;48m \033[48;2;101;65;52m \033[48;2;102;66;52m \033[48;2;97;61;48m \033[48;2;94;58;43m \033[48;2;89;53;38m \033[48;2;94;58;42m \033[48;2;92;57;45m \033[48;2;90;55;43m \033[48;2;94;59;47m \033[48;2;104;67;59m \033[48;2;103;67;58m \033[48;2;103;66;58m \033[48;2;105;67;58m \033[48;2;115;79;70m \033[48;2;117;80;71m \033[48;2;115;85;77m \033[48;2;147;121;115m \033[48;2;186;163;173m \033[48;2;178;162;177m \033[48;2;176;156;180m \033[48;2;176;156;183m \033[48;2;176;159;185m \033[48;2;175;159;185m \033[48;2;174;158;184m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;173;159;185m \033[48;2;170;156;182m \033[48;2;168;154;180m \033[48;2;173;159;185m \033[48;2;167;153;179m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;149;175m \033[48;2;166;152;178m \033[48;2;172;158;184m \033[48;2;174;160;186m \033[48;2;174;160;186m \033[48;2;176;162;188m \033[48;2;173;157;184m \033[48;2;172;156;183m \033[48;2;172;156;183m \033[48;2;165;148;178m \033[48;2;165;148;180m \033[48;2;164;151;181m \033[48;2;162;152;179m \033[48;2;162;152;177m \033[48;2;162;152;178m \033[48;2;162;152;179m \033[48;2;162;151;181m \033[48;2;163;152;182m \033[m");
$display("\033[48;2;183;172;204m \033[48;2;183;172;204m \033[48;2;185;172;202m \033[48;2;181;168;198m \033[48;2;178;165;195m \033[48;2;180;167;197m \033[48;2;187;174;204m \033[48;2;183;170;200m \033[48;2;180;167;197m \033[48;2;179;166;196m \033[48;2;172;159;190m \033[48;2;172;159;185m \033[48;2;172;159;185m \033[48;2;176;163;189m \033[48;2;181;167;192m \033[48;2;184;170;195m \033[48;2;184;170;195m \033[48;2;183;169;195m \033[48;2;181;167;193m \033[48;2;170;156;182m \033[48;2;172;156;183m \033[48;2;171;155;182m \033[48;2;170;154;181m \033[48;2;170;154;181m \033[48;2;166;150;178m \033[48;2;166;150;177m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;148;174m \033[48;2;164;149;172m \033[48;2;164;149;170m \033[48;2;165;151;168m \033[48;2;166;145;163m \033[48;2;177;146;147m \033[48;2;189;145;128m \033[48;2;196;140;109m \033[48;2;166;97;69m \033[48;2;157;82;49m \033[48;2;168;99;71m \033[48;2;173;109;81m \033[48;2;150;92;65m \033[48;2;142;85;64m \033[48;2;143;85;70m \033[48;2;144;92;80m \033[48;2;143;91;87m \033[48;2;141;92;88m \033[48;2;138;90;90m \033[48;2;140;92;90m \033[48;2;142;93;96m \033[48;2;152;102;113m \033[48;2;148;108;108m \033[48;2;148;108;108m \033[48;2;151;111;112m \033[48;2;147;108;113m \033[48;2;141;102;106m \033[48;2;137;98;103m \033[48;2;138;98;105m \033[48;2;148;108;118m \033[48;2;149;110;118m \033[48;2;154;114;119m \033[48;2;154;115;120m \033[48;2;153;114;118m \033[48;2;146;109;103m \033[48;2;142;105;99m \033[48;2;130;93;88m \033[48;2;116;79;70m \033[48;2;102;65;58m \033[48;2;107;70;62m \033[48;2;102;65;56m \033[48;2;108;71;62m \033[48;2;111;74;65m \033[48;2;116;83;78m \033[48;2;132;108;98m \033[48;2;176;155;152m \033[48;2;178;160;175m \033[48;2;176;156;181m \033[48;2;176;156;183m \033[48;2;176;159;185m \033[48;2;175;159;185m \033[48;2;174;158;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;173;159;185m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;175;161;187m \033[48;2;173;159;185m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;149;175m \033[48;2;166;152;178m \033[48;2;172;158;184m \033[48;2;175;161;187m \033[48;2;175;161;187m \033[48;2;177;163;189m \033[48;2;176;159;186m \033[48;2;174;158;185m \033[48;2;175;159;186m \033[48;2;170;151;182m \033[48;2;166;149;181m \033[48;2;164;151;181m \033[48;2;162;152;179m \033[48;2;162;152;177m \033[48;2;162;152;177m \033[48;2;162;152;177m \033[48;2;163;153;177m \033[48;2;163;153;177m \033[m");
$display("\033[48;2;180;169;201m \033[48;2;177;166;198m \033[48;2;176;165;195m \033[48;2;179;168;198m \033[48;2;177;166;196m \033[48;2;181;170;202m \033[48;2;180;169;201m \033[48;2;184;173;205m \033[48;2;187;174;204m \033[48;2;183;170;200m \033[48;2;179;166;196m \033[48;2;182;169;195m \033[48;2;184;171;197m \033[48;2;181;168;194m \033[48;2;189;177;201m \033[48;2;190;176;201m \033[48;2;189;173;199m \033[48;2;189;173;200m \033[48;2;190;174;201m \033[48;2;184;168;195m \033[48;2;177;161;188m \033[48;2;176;160;187m \033[48;2;170;154;181m \033[48;2;171;155;181m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;148;174m \033[48;2;167;147;172m \033[48;2;167;148;169m \033[48;2;168;149;168m \033[48;2;170;145;159m \033[48;2;181;144;145m \033[48;2;192;143;129m \033[48;2;194;134;105m \033[48;2;160;95;61m \033[48;2;132;66;37m \033[48;2;118;60;39m \033[48;2;117;70;51m \033[48;2;134;89;73m \033[48;2;141;93;78m \033[48;2;146;97;86m \033[48;2;143;94;91m \033[48;2;139;87;91m \033[48;2;136;84;88m \033[48;2;136;84;88m \033[48;2;142;86;93m \033[48;2;148;92;101m \033[48;2;153;102;111m \033[48;2;152;104;116m \033[48;2;155;107;119m \033[48;2;158;110;122m \033[48;2;157;114;123m \033[48;2;157;114;123m \033[48;2;158;115;124m \033[48;2;160;117;128m \033[48;2;159;113;128m \033[48;2;161;117;134m \033[48;2;160;114;139m \033[48;2;160;114;136m \033[48;2;163;117;137m \033[48;2;164;119;132m \033[48;2;162;117;131m \033[48;2;162;116;132m \033[48;2;160;114;126m \033[48;2;148;103;109m \033[48;2;119;76;75m \033[48;2;107;68;61m \033[48;2;105;68;61m \033[48;2;102;68;59m \033[48;2;105;76;63m \033[48;2;131;106;100m \033[48;2;175;154;155m \033[48;2;172;158;174m \033[48;2;170;155;174m \033[48;2;169;154;176m \033[48;2;173;157;183m \033[48;2;173;157;183m \033[48;2;174;158;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;172;158;184m \033[48;2;174;160;186m \033[48;2;172;158;184m \033[48;2;169;155;181m \033[48;2;172;158;184m \033[48;2;172;158;184m \033[48;2;167;153;179m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;165;148;174m \033[48;2;166;151;177m \033[48;2;168;156;182m \033[48;2;171;159;185m \033[48;2;171;158;184m \033[48;2;168;155;181m \033[48;2;168;155;182m \033[48;2;166;153;183m \033[48;2;171;158;188m \033[48;2;172;159;189m \033[48;2;170;159;187m \033[48;2;167;155;185m \033[48;2;163;151;181m \033[48;2;162;151;181m \033[48;2;162;151;181m \033[48;2;162;151;181m \033[48;2;162;152;179m \033[48;2;163;153;180m \033[m");
$display("\033[48;2;178;167;197m \033[48;2;185;174;204m \033[48;2;187;177;202m \033[48;2;185;175;200m \033[48;2;185;175;200m \033[48;2;184;173;203m \033[48;2;179;168;198m \033[48;2;178;167;197m \033[48;2;182;171;201m \033[48;2;183;172;202m \033[48;2;177;166;197m \033[48;2;181;171;196m \033[48;2;184;174;199m \033[48;2;181;171;196m \033[48;2;182;169;195m \033[48;2;185;171;197m \033[48;2;186;170;197m \033[48;2;186;172;197m \033[48;2;186;172;197m \033[48;2;186;172;197m \033[48;2;185;169;195m \033[48;2;182;166;192m \033[48;2;182;166;192m \033[48;2;189;169;196m \033[48;2;182;161;189m \033[48;2;174;154;181m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;149;171m \033[48;2;168;149;168m \033[48;2;170;147;165m \033[48;2;177;146;153m \033[48;2;186;145;143m \033[48;2;193;139;126m \033[48;2;168;101;79m \033[48;2;121;50;28m \033[48;2;119;53;37m \033[48;2;116;66;48m \033[48;2;118;80;67m \033[48;2;130;93;90m \033[48;2;140;91;94m \033[48;2;142;93;96m \033[48;2;138;89;92m \033[48;2;137;84;89m \033[48;2;137;85;89m \033[48;2;137;85;89m \033[48;2;139;88;90m \033[48;2;144;94;97m \033[48;2;148;97;104m \033[48;2;145;100;105m \033[48;2;150;103;111m \033[48;2;153;105;117m \033[48;2;155;107;121m \033[48;2;155;107;121m \033[48;2;156;108;122m \033[48;2;159;110;129m \033[48;2;159;110;131m \033[48;2;160;110;134m \033[48;2;161;111;136m \033[48;2;161;111;136m \033[48;2;163;113;138m \033[48;2;164;114;141m \033[48;2;167;117;144m \033[48;2;163;113;140m \033[48;2;162;112;135m \033[48;2;159;110;130m \033[48;2;146;99;109m \033[48;2;112;72;73m \033[48;2;103;66;61m \033[48;2;101;68;57m \033[48;2;109;79;68m \033[48;2;141;118;112m \033[48;2;181;162;167m \033[48;2;174;156;174m \033[48;2;174;155;175m \033[48;2;175;156;179m \033[48;2;181;161;188m \033[48;2;181;161;188m \033[48;2;179;159;186m \033[48;2;179;161;189m \033[48;2;175;159;186m \033[48;2;172;156;183m \033[48;2;172;158;184m \033[48;2;172;158;184m \033[48;2;168;154;180m \033[48;2;167;153;179m \033[48;2;169;155;181m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;148;178m \033[48;2;166;152;182m \033[48;2;169;157;188m \033[48;2;172;161;191m \033[48;2;172;161;192m \033[48;2;172;161;191m \033[48;2;171;160;190m \033[48;2;171;160;190m \033[48;2;173;164;194m \033[48;2;174;163;193m \033[48;2;170;159;189m \033[48;2;166;155;185m \033[48;2;162;151;181m \033[48;2;162;151;181m \033[48;2;162;151;181m \033[48;2;162;151;181m \033[48;2;161;150;180m \033[48;2;162;151;181m \033[m");
$display("\033[48;2;183;172;202m \033[48;2;179;168;198m \033[48;2;183;173;198m \033[48;2;186;176;201m \033[48;2;186;176;201m \033[48;2;187;177;206m \033[48;2;188;177;207m \033[48;2;182;171;201m \033[48;2;181;170;200m \033[48;2;178;168;197m \033[48;2;180;169;199m \033[48;2;178;167;193m \033[48;2;178;169;193m \033[48;2;179;170;195m \033[48;2;179;167;196m \033[48;2;177;163;189m \033[48;2;178;161;189m \033[48;2;175;161;186m \033[48;2;171;157;182m \033[48;2;170;156;181m \033[48;2;172;156;182m \033[48;2;176;160;186m \033[48;2;174;158;184m \033[48;2;182;162;189m \033[48;2;183;163;190m \033[48;2;183;163;190m \033[48;2;173;153;178m \033[48;2;168;148;173m \033[48;2;167;147;172m \033[48;2;166;148;170m \033[48;2;167;148;168m \033[48;2;170;147;165m \033[48;2;181;147;150m \033[48;2;192;146;140m \033[48;2;189;130;111m \033[48;2;153;81;63m \033[48;2;124;58;33m \033[48;2;118;70;48m \033[48;2;117;77;55m \033[48;2;123;85;73m \033[48;2;135;90;90m \033[48;2;140;91;94m \033[48;2;141;91;94m \033[48;2;137;88;91m \033[48;2;133;87;89m \033[48;2;133;87;89m \033[48;2;135;87;90m \033[48;2;133;89;88m \033[48;2;136;92;93m \033[48;2;139;94;99m \033[48;2;145;98;104m \033[48;2;148;101;109m \033[48;2;153;105;117m \033[48;2;156;108;123m \033[48;2;159;111;125m \033[48;2;160;112;126m \033[48;2;157;107;127m \033[48;2;159;110;131m \033[48;2;158;109;133m \033[48;2;160;110;135m \033[48;2;163;113;138m \033[48;2;163;113;138m \033[48;2;165;115;142m \033[48;2;165;115;142m \033[48;2;163;113;140m \033[48;2;162;112;134m \033[48;2;159;110;129m \033[48;2;153;105;115m \033[48;2;127;85;86m \033[48;2;121;83;80m \033[48;2;109;75;67m \033[48;2;120;89;82m \033[48;2;165;141;140m \033[48;2;178;159;171m \033[48;2;170;151;170m \033[48;2;170;151;171m \033[48;2;174;155;177m \033[48;2;179;159;186m \033[48;2;179;159;186m \033[48;2;179;159;186m \033[48;2;178;159;187m \033[48;2;176;160;187m \033[48;2;173;157;184m \033[48;2;176;162;188m \033[48;2;176;162;188m \033[48;2;172;159;184m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;148;178m \033[48;2;166;152;182m \033[48;2;168;156;186m \033[48;2;171;160;190m \033[48;2;171;160;190m \033[48;2;175;164;194m \033[48;2;173;162;192m \033[48;2;173;162;192m \033[48;2;172;162;192m \033[48;2;165;154;184m \033[48;2;163;152;182m \033[48;2;161;151;181m \033[48;2;160;149;179m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;162;151;181m \033[m");
$display("\033[48;2;187;177;202m \033[48;2;185;175;200m \033[48;2;183;173;198m \033[48;2;184;174;199m \033[48;2;180;170;195m \033[48;2;178;168;193m \033[48;2;174;164;189m \033[48;2;174;164;189m \033[48;2;175;161;194m \033[48;2;173;159;192m \033[48;2;174;160;193m \033[48;2;178;163;197m \033[48;2;181;168;197m \033[48;2;185;172;198m \033[48;2;190;176;201m \033[48;2;186;172;197m \033[48;2;184;170;195m \033[48;2;192;178;203m \033[48;2;191;177;202m \033[48;2;189;175;200m \033[48;2;190;174;200m \033[48;2;189;173;199m \033[48;2;183;167;193m \033[48;2;190;170;197m \033[48;2;185;165;192m \033[48;2;174;154;181m \033[48;2;171;151;176m \033[48;2;169;149;174m \033[48;2;168;148;173m \033[48;2;167;149;171m \033[48;2;168;149;169m \033[48;2;170;147;165m \033[48;2;179;145;146m \033[48;2;186;139;124m \033[48;2;160;98;78m \033[48;2;145;80;53m \033[48;2;122;67;41m \033[48;2;114;72;50m \033[48;2;123;87;71m \033[48;2;131;93;83m \033[48;2;139;98;95m \033[48;2;136;90;92m \033[48;2;135;89;91m \033[48;2;127;80;82m \033[48;2;130;82;80m \033[48;2;129;81;79m \033[48;2;130;82;80m \033[48;2;133;87;87m \033[48;2;133;87;89m \033[48;2;131;84;90m \033[48;2;140;93;99m \033[48;2;149;102;110m \033[48;2;156;107;119m \033[48;2;155;105;125m \033[48;2;162;113;131m \033[48;2;158;109;128m \033[48;2;154;106;119m \033[48;2;157;109;123m \033[48;2;158;109;128m \033[48;2;161;111;134m \033[48;2;164;114;139m \033[48;2;165;115;140m \033[48;2;165;115;140m \033[48;2;162;112;137m \033[48;2;164;114;139m \033[48;2;164;115;137m \033[48;2;161;114;130m \033[48;2;149;101;114m \033[48;2;130;89;92m \033[48;2;120;81;82m \033[48;2;111;76;72m \033[48;2;111;85;78m \033[48;2;164;142;144m \033[48;2;173;156;168m \033[48;2;172;153;172m \033[48;2;172;153;173m \033[48;2;175;156;179m \033[48;2;177;157;182m \033[48;2;181;161;186m \033[48;2;179;159;184m \033[48;2;178;159;187m \033[48;2;176;160;187m \033[48;2;174;158;185m \033[48;2;179;163;190m \033[48;2;179;163;190m \033[48;2;178;162;189m \033[48;2;170;157;182m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;162;148;178m \033[48;2;165;151;181m \033[48;2;168;156;187m \033[48;2;168;158;185m \033[48;2;172;162;187m \033[48;2;172;162;187m \033[48;2;172;161;189m \033[48;2;172;159;189m \033[48;2;167;154;184m \033[48;2;164;151;181m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;162;150;180m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;161;150;180m \033[48;2;162;151;181m \033[m");
$display("\033[48;2;183;173;198m \033[48;2;186;176;202m \033[48;2;187;177;202m \033[48;2;187;177;202m \033[48;2;190;180;205m \033[48;2;191;181;206m \033[48;2;189;179;204m \033[48;2;189;179;204m \033[48;2;189;176;207m \033[48;2;180;166;197m \033[48;2;180;165;197m \033[48;2;186;173;203m \033[48;2;187;172;203m \033[48;2;190;172;205m \033[48;2;188;173;204m \033[48;2;184;169;200m \033[48;2;183;168;199m \033[48;2;190;176;202m \033[48;2;191;177;203m \033[48;2;189;175;201m \033[48;2;190;174;200m \033[48;2;187;171;197m \033[48;2;183;167;193m \033[48;2;175;159;185m \033[48;2;171;155;181m \033[48;2;169;153;179m \033[48;2;168;152;179m \033[48;2;166;150;176m \033[48;2;165;150;173m \033[48;2;170;148;171m \033[48;2;171;147;169m \033[48;2;171;146;165m \033[48;2;177;141;141m \033[48;2;177;128;110m \033[48;2;175;120;88m \033[48;2;153;98;70m \033[48;2;126;76;51m \033[48;2;127;85;65m \033[48;2;137;92;85m \033[48;2;141;96;91m \033[48;2;137;91;88m \033[48;2;136;86;89m \033[48;2;130;80;83m \033[48;2;129;79;84m \033[48;2;127;77;76m \033[48;2;129;82;79m \033[48;2;127;83;80m \033[48;2;129;79;83m \033[48;2;123;74;78m \033[48;2;114;65;69m \033[48;2;116;65;70m \033[48;2;118;67;72m \033[48;2;130;79;83m \033[48;2;136;85;92m \033[48;2;153;102;109m \033[48;2;155;104;111m \033[48;2;144;95;108m \033[48;2;145;95;108m \033[48;2;153;103;114m \033[48;2;158;111;130m \033[48;2;164;118;136m \033[48;2;164;114;139m \033[48;2;166;115;141m \033[48;2;166;117;139m \033[48;2;159;110;130m \033[48;2;158;110;126m \033[48;2;161;113;127m \033[48;2;149;102;113m \033[48;2;128;84;86m \033[48;2;117;77;77m \033[48;2;110;78;73m \033[48;2;130;112;103m \033[48;2;172;153;153m \033[48;2;171;154;169m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;169;149;174m \033[48;2;171;151;178m \033[48;2;174;154;181m \033[48;2;174;154;181m \033[48;2;174;154;185m \033[48;2;172;155;187m \033[48;2;170;153;185m \033[48;2;177;161;189m \033[48;2;177;161;188m \033[48;2;177;161;188m \033[48;2;173;157;184m \033[48;2;167;151;178m \033[48;2;166;150;177m \033[48;2;165;149;179m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;165;150;181m \033[48;2;164;149;180m \033[48;2;172;157;188m \033[48;2;175;162;192m \033[48;2;173;162;192m \033[48;2;178;167;197m \033[48;2;177;164;194m \033[48;2;173;158;189m \033[48;2;172;157;188m \033[48;2;167;152;183m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[48;2;164;150;180m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;161;150;180m \033[48;2;162;151;181m \033[m");
$display("\033[48;2;189;178;210m \033[48;2;192;181;214m \033[48;2;187;177;202m \033[48;2;186;176;203m \033[48;2;189;179;205m \033[48;2;189;179;204m \033[48;2;188;178;205m \033[48;2;188;178;204m \033[48;2;189;176;202m \033[48;2;179;166;192m \033[48;2;184;171;198m \033[48;2;187;174;204m \033[48;2;187;172;202m \033[48;2;187;171;201m \033[48;2;187;172;203m \033[48;2;182;167;198m \033[48;2;185;170;201m \033[48;2;190;176;202m \033[48;2;187;173;199m \033[48;2;177;163;189m \033[48;2;175;157;183m \033[48;2;173;156;181m \033[48;2;170;154;180m \033[48;2;172;155;181m \033[48;2;172;155;181m \033[48;2;172;154;181m \033[48;2;168;152;179m \033[48;2;166;150;176m \033[48;2;165;150;173m \033[48;2;170;148;171m \033[48;2;171;147;169m \033[48;2;173;146;165m \033[48;2;172;141;145m \033[48;2;175;132;119m \033[48;2;156;106;82m \033[48;2;134;80;54m \033[48;2;143;92;68m \033[48;2;131;90;69m \033[48;2;138;94;87m \033[48;2;137;91;86m \033[48;2;136;91;89m \033[48;2;137;87;90m \033[48;2;137;88;91m \033[48;2;120;71;74m \033[48;2;114;64;63m \033[48;2;105;58;55m \033[48;2;96;53;50m \033[48;2;105;58;62m \033[48;2;121;74;77m \033[48;2;116;69;74m \033[48;2;123;72;78m \033[48;2;125;75;79m \033[48;2;118;67;72m \033[48;2;125;74;80m \033[48;2;145;94;102m \033[48;2;162;111;118m \033[48;2;150;94;103m \033[48;2;134;78;87m \033[48;2;125;68;77m \033[48;2;119;67;71m \033[48;2;117;65;73m \033[48;2;124;72;82m \033[48;2;131;83;99m \033[48;2;135;87;102m \033[48;2;152;104;116m \033[48;2;160;112;128m \033[48;2;152;104;117m \033[48;2;146;98;108m \033[48;2;117;72;76m \033[48;2;113;75;74m \033[48;2;117;87;81m \033[48;2;141;122;118m \033[48;2;176;157;162m \033[48;2;170;152;172m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;168;148;173m \033[48;2;170;150;177m \033[48;2;166;146;173m \033[48;2;170;150;177m \033[48;2;175;156;187m \033[48;2;173;156;188m \033[48;2;178;161;193m \033[48;2;181;165;195m \033[48;2;178;162;189m \033[48;2;179;163;190m \033[48;2;173;157;184m \033[48;2;170;154;181m \033[48;2;165;149;176m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;170;155;186m \033[48;2;177;164;194m \033[48;2;175;164;194m \033[48;2;177;166;196m \033[48;2;179;165;196m \033[48;2;176;161;192m \033[48;2;178;163;194m \033[48;2;176;162;192m \033[48;2;168;152;184m \033[48;2;167;152;183m \033[48;2;164;151;181m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;161;150;180m \033[48;2;162;151;181m \033[m");
$display("\033[48;2;174;163;197m \033[48;2;177;166;200m \033[48;2;181;170;200m \033[48;2;186;175;205m \033[48;2;190;179;209m \033[48;2;188;177;207m \033[48;2;185;174;204m \033[48;2;188;177;207m \033[48;2;185;172;198m \033[48;2;181;168;194m \033[48;2;187;174;200m \033[48;2;188;174;200m \033[48;2;188;174;200m \033[48;2;188;174;200m \033[48;2;187;172;203m \033[48;2;184;169;200m \033[48;2;191;176;207m \033[48;2;190;176;202m \033[48;2;178;164;190m \033[48;2;172;158;184m \033[48;2;177;157;184m \033[48;2;177;157;184m \033[48;2;177;157;184m \033[48;2;175;155;182m \033[48;2;175;155;182m \033[48;2;172;151;179m \033[48;2;167;151;177m \033[48;2;167;151;177m \033[48;2;164;148;174m \033[48;2;167;148;170m \033[48;2;170;146;167m \033[48;2;189;147;172m \033[48;2;186;136;142m \033[48;2;183;129;124m \033[48;2;169;115;101m \033[48;2;181;126;103m \033[48;2;178;128;101m \033[48;2;184;142;121m \033[48;2;185;139;124m \033[48;2;171;124;116m \033[48;2;144;97;95m \033[48;2;137;88;91m \033[48;2;136;87;90m \033[48;2;138;89;92m \033[48;2;138;93;94m \033[48;2;140;96;97m \033[48;2;140;100;100m \033[48;2;143;103;103m \033[48;2;143;102;106m \033[48;2;135;87;96m \033[48;2;128;78;88m \033[48;2;123;74;80m \033[48;2;127;78;82m \033[48;2;133;83;84m \033[48;2;147;98;100m \033[48;2;159;108;115m \033[48;2;165;114;126m \033[48;2;159;107;119m \033[48;2;124;73;84m \033[48;2;114;61;69m \033[48;2;103;50;57m \033[48;2;117;71;76m \033[48;2;144;95;106m \033[48;2;155;107;119m \033[48;2;149;101;113m \033[48;2;144;96;111m \033[48;2;147;99;112m \033[48;2;146;99;108m \033[48;2;109;71;70m \033[48;2;115;83;80m \033[48;2;141;121;114m \033[48;2;180;164;166m \033[48;2;172;154;170m \033[48;2;169;150;170m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;167;147;174m \033[48;2;167;147;174m \033[48;2;167;147;174m \033[48;2;168;148;175m \033[48;2;167;148;178m \033[48;2;165;148;180m \033[48;2;168;151;183m \033[48;2;175;159;187m \033[48;2;178;162;189m \033[48;2;178;162;189m \033[48;2;179;163;190m \033[48;2;171;155;182m \033[48;2;166;150;177m \033[48;2;165;149;179m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;168;153;184m \033[48;2;175;162;192m \033[48;2;173;162;192m \033[48;2;175;164;194m \033[48;2;177;164;194m \033[48;2;172;159;189m \033[48;2;172;159;189m \033[48;2;166;153;183m \033[48;2;165;152;182m \033[48;2;164;151;181m \033[48;2;164;151;180m \033[48;2;164;151;179m \033[48;2;164;151;179m \033[48;2;164;151;179m \033[48;2;164;151;181m \033[48;2;164;151;181m \033[m");
$display("\033[48;2;175;164;198m \033[48;2;175;164;198m \033[48;2;175;164;194m \033[48;2;182;171;201m \033[48;2;189;178;208m \033[48;2;186;175;205m \033[48;2;184;173;203m \033[48;2;185;174;204m \033[48;2;181;168;198m \033[48;2;180;167;197m \033[48;2;183;170;201m \033[48;2;182;168;194m \033[48;2;179;165;191m \033[48;2;182;167;193m \033[48;2;183;167;194m \033[48;2;183;167;194m \033[48;2;185;169;196m \033[48;2;183;166;198m \033[48;2;176;159;191m \033[48;2;174;157;189m \033[48;2;174;154;181m \033[48;2;174;154;181m \033[48;2;174;154;181m \033[48;2;173;153;180m \033[48;2;173;153;180m \033[48;2;172;152;179m \033[48;2;171;151;176m \033[48;2;169;149;174m \033[48;2;167;147;172m \033[48;2;173;141;166m \033[48;2;176;116;143m \033[48;2;170;60;92m \033[48;2;189;57;88m \033[48;2;190;64;86m \033[48;2;173;74;76m \033[48;2;185;116;100m \033[48;2;206;156;134m \033[48;2;187;142;117m \033[48;2;188;139;125m \033[48;2;178;123;113m \033[48;2;154;105;98m \033[48;2;140;91;87m \033[48;2;136;88;85m \033[48;2;138;95;96m \033[48;2;146;101;106m \033[48;2;146;100;106m \033[48;2;146;102;107m \033[48;2;146;99;105m \033[48;2;136;88;94m \033[48;2;127;80;86m \033[48;2;124;75;79m \033[48;2;127;78;81m \033[48;2;132;84;81m \033[48;2;137;89;90m \033[48;2;148;99;104m \033[48;2;159;109;118m \033[48;2;160;112;128m \033[48;2;160;111;130m \033[48;2;156;107;129m \033[48;2;150;102;124m \033[48;2;150;101;124m \033[48;2;158;109;133m \033[48;2;157;108;129m \033[48;2;140;91;112m \033[48;2;145;96;116m \033[48;2;154;105;125m \033[48;2;156;108;124m \033[48;2;135;93;105m \033[48;2;131;101;97m \033[48;2;183;157;159m \033[48;2;172;152;161m \033[48;2;170;154;175m \033[48;2;166;151;171m \033[48;2;166;151;171m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;168;148;175m \033[48;2;165;147;178m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;170;153;185m \033[48;2;174;158;187m \033[48;2;172;156;183m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;165;151;177m \033[48;2;169;155;181m \033[48;2;169;156;182m \033[48;2;167;154;181m \033[48;2;165;152;181m \033[48;2;163;150;180m \033[48;2;164;151;181m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;164;151;181m \033[48;2;165;150;179m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;165;151;179m \033[48;2;165;150;181m \033[48;2;165;150;181m \033[m");
$display("\033[48;2;173;162;196m \033[48;2;173;162;196m \033[48;2;174;163;195m \033[48;2;185;175;204m \033[48;2;190;180;207m \033[48;2;189;179;205m \033[48;2;188;179;206m \033[48;2;188;178;204m \033[48;2;181;168;198m \033[48;2;183;170;200m \033[48;2;188;175;205m \033[48;2;189;175;201m \033[48;2;187;173;199m \033[48;2;188;174;200m \033[48;2;183;168;195m \033[48;2;175;160;186m \033[48;2;174;159;186m \033[48;2;173;156;188m \033[48;2;174;157;189m \033[48;2;173;156;188m \033[48;2;174;154;181m \033[48;2;174;154;181m \033[48;2;174;154;181m \033[48;2;173;153;179m \033[48;2;171;151;177m \033[48;2;171;151;176m \033[48;2;169;150;173m \033[48;2;169;149;173m \033[48;2;169;149;173m \033[48;2;174;135;162m \033[48;2;169;102;135m \033[48;2;169;61;92m \033[48;2;185;50;88m \033[48;2;191;48;83m \033[48;2;179;64;84m \033[48;2;166;90;87m \033[48;2;196;142;131m \033[48;2;177;127;113m \033[48;2;171;117;104m \033[48;2;155;98;91m \033[48;2;146;90;87m \033[48;2;140;91;88m \033[48;2;138;89;87m \033[48;2;135;88;87m \033[48;2;138;88;93m \033[48;2;138;88;93m \033[48;2;137;85;92m \033[48;2;133;82;87m \033[48;2;129;78;84m \033[48;2;127;76;82m \033[48;2;131;80;84m \033[48;2;130;80;83m \033[48;2;136;85;90m \033[48;2;143;93;100m \033[48;2;158;107;120m \033[48;2;163;110;124m \033[48;2;161;111;126m \033[48;2;164;114;132m \033[48;2;169;118;138m \033[48;2;164;116;137m \033[48;2;161;111;138m \033[48;2;160;110;138m \033[48;2;162;112;138m \033[48;2;165;115;140m \033[48;2;163;114;137m \033[48;2;160;113;134m \033[48;2;159;113;129m \033[48;2;130;91;103m \033[48;2;166;139;145m \033[48;2;179;157;168m \033[48;2;175;160;176m \033[48;2;171;153;178m \033[48;2;168;149;174m \033[48;2;168;150;175m \033[48;2;168;148;174m \033[48;2;168;148;174m \033[48;2;168;148;174m \033[48;2;168;148;174m \033[48;2;168;148;174m \033[48;2;168;148;174m \033[48;2;167;148;177m \033[48;2;165;149;178m \033[48;2;165;148;177m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;167;150;180m \033[48;2;169;153;182m \033[48;2;167;150;179m \033[48;2;165;149;179m \033[48;2;165;149;178m \033[48;2;165;149;178m \033[48;2;164;149;178m \033[48;2;164;149;178m \033[48;2;167;152;181m \033[48;2;173;159;186m \033[48;2;173;159;185m \033[48;2;165;151;177m \033[48;2;164;151;180m \033[48;2;164;151;181m \033[48;2;164;151;181m \033[48;2;164;150;180m \033[48;2;164;150;180m \033[48;2;163;151;181m \033[48;2;163;150;179m \033[48;2;164;151;177m \033[48;2;165;151;177m \033[48;2;165;151;180m \033[48;2;169;155;185m \033[48;2;167;154;184m \033[m");
$display("\033[48;2;172;161;195m \033[48;2;175;164;198m \033[48;2;175;164;196m \033[48;2;182;172;198m \033[48;2;187;177;202m \033[48;2;187;177;202m \033[48;2;189;179;204m \033[48;2;186;176;201m \033[48;2;178;165;195m \033[48;2;184;171;201m \033[48;2;188;174;205m \033[48;2;178;164;190m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;172;155;187m \033[48;2;172;155;187m \033[48;2;171;154;186m \033[48;2;174;154;181m \033[48;2;171;151;178m \033[48;2;172;152;179m \033[48;2;172;152;177m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;170;151;173m \033[48;2;170;151;173m \033[48;2;169;150;172m \033[48;2;177;147;171m \033[48;2;183;139;164m \033[48;2;175;94;119m \033[48;2;168;51;83m \033[48;2;195;54;91m \033[48;2;184;60;90m \033[48;2;167;73;89m \033[48;2;165;101;104m \033[48;2;175;124;120m \033[48;2;158;109;102m \033[48;2;146;97;92m \033[48;2;139;89;87m \033[48;2;137;87;86m \033[48;2;136;86;85m \033[48;2;135;85;84m \033[48;2;135;82;88m \033[48;2;132;79;85m \033[48;2;133;80;86m \033[48;2;135;79;85m \033[48;2;131;75;82m \033[48;2;124;69;74m \033[48;2;125;67;73m \033[48;2;105;47;53m \033[48;2;117;61;66m \033[48;2;123;68;74m \033[48;2;133;75;84m \033[48;2;146;90;103m \033[48;2;152;102;114m \033[48;2;159;108;126m \033[48;2;163;112;131m \033[48;2;165;116;138m \033[48;2;168;118;145m \033[48;2;169;119;148m \033[48;2;166;116;143m \033[48;2;163;112;138m \033[48;2;162;113;135m \033[48;2;161;109;131m \033[48;2;157;109;125m \033[48;2;142;97;111m \033[48;2;140;98;114m \033[48;2;185;152;169m \033[48;2;179;151;173m \033[48;2;178;158;183m \033[48;2;175;155;180m \033[48;2;171;151;176m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;148;176m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;164;147;179m \033[48;2;165;148;180m \033[48;2;165;148;180m \033[48;2;165;148;180m \033[48;2;165;148;180m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;165;150;181m \033[48;2;167;152;180m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;151;180m \033[48;2;164;151;181m \033[48;2;164;151;181m \033[48;2;164;149;180m \033[48;2;164;149;180m \033[48;2;162;151;181m \033[48;2;162;151;178m \033[48;2;163;150;176m \033[48;2;162;149;175m \033[48;2;165;152;180m \033[48;2;170;157;187m \033[48;2;172;159;189m \033[m");
$display("\033[48;2;175;164;198m \033[48;2;175;164;198m \033[48;2;175;164;194m \033[48;2;173;162;192m \033[48;2;180;169;199m \033[48;2;187;174;204m \033[48;2;192;179;209m \033[48;2;188;175;205m \033[48;2;182;169;199m \033[48;2;182;169;199m \033[48;2;175;162;192m \033[48;2;172;157;188m \033[48;2;170;155;186m \033[48;2;170;155;186m \033[48;2;170;155;186m \033[48;2;171;156;187m \033[48;2;171;156;187m \033[48;2;171;154;186m \033[48;2;171;154;186m \033[48;2;171;154;186m \033[48;2;171;155;181m \033[48;2;171;155;181m \033[48;2;171;155;181m \033[48;2;174;154;179m \033[48;2;173;153;178m \033[48;2;173;153;178m \033[48;2;173;154;176m \033[48;2;173;154;176m \033[48;2;174;155;177m \033[48;2;176;154;175m \033[48;2;181;149;167m \033[48;2;176;128;147m \033[48;2;157;96;111m \033[48;2;154;87;104m \033[48;2;140;79;90m \033[48;2;150;82;87m \033[48;2;142;82;83m \033[48;2;152;103;101m \033[48;2;154;104;103m \033[48;2;148;98;97m \033[48;2;145;95;94m \033[48;2;142;92;95m \033[48;2;138;88;91m \033[48;2;136;86;89m \033[48;2;135;83;87m \033[48;2;135;83;87m \033[48;2;134;82;86m \033[48;2;131;79;81m \033[48;2;129;77;81m \033[48;2;127;74;82m \033[48;2;133;76;85m \033[48;2;136;79;88m \033[48;2;144;87;96m \033[48;2;153;97;110m \033[48;2;156;100;113m \033[48;2;155;100;112m \033[48;2;154;102;119m \033[48;2;166;115;133m \033[48;2;152;100;123m \033[48;2;156;107;129m \033[48;2;159;110;132m \033[48;2;161;112;134m \033[48;2;160;111;132m \033[48;2;157;108;127m \033[48;2;157;109;124m \033[48;2;158;110;126m \033[48;2;157;107;124m \033[48;2;165;111;129m \033[48;2;146;88;108m \033[48;2;186;140;161m \033[48;2;183;154;176m \033[48;2;178;157;183m \033[48;2;177;157;182m \033[48;2;175;155;180m \033[48;2;176;159;182m \033[48;2;172;157;180m \033[48;2;166;151;174m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;174m \033[48;2;164;148;175m \033[48;2;164;148;175m \033[48;2;164;148;175m \033[48;2;163;149;175m \033[48;2;163;149;175m \033[48;2;163;149;175m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;163;150;178m \033[48;2;163;150;180m \033[48;2;163;150;180m \033[48;2;164;150;179m \033[48;2;165;151;177m \033[48;2;170;156;182m \033[48;2;176;162;189m \033[48;2;175;160;191m \033[48;2;176;161;192m \033[m");
$display("\033[48;2;175;164;196m \033[48;2;175;164;196m \033[48;2;177;163;196m \033[48;2;175;161;194m \033[48;2;175;161;194m \033[48;2;178;165;195m \033[48;2;184;171;201m \033[48;2;183;170;200m \033[48;2;177;162;193m \033[48;2;174;159;190m \033[48;2;174;159;190m \033[48;2;172;157;188m \033[48;2;170;155;186m \033[48;2;171;156;187m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;171;155;181m \033[48;2;169;153;179m \033[48;2;168;152;178m \033[48;2;173;153;178m \033[48;2;174;154;179m \033[48;2;179;159;184m \033[48;2;178;159;181m \033[48;2;175;156;178m \033[48;2;174;155;177m \033[48;2;171;152;171m \033[48;2;172;153;171m \033[48;2;171;153;171m \033[48;2;179;150;165m \033[48;2;159;113;128m \033[48;2;152;87;100m \033[48;2;150;82;91m \033[48;2;146;87;89m \033[48;2;142;93;85m \033[48;2;148;100;98m \033[48;2;145;97;95m \033[48;2;142;94;92m \033[48;2;141;91;94m \033[48;2;141;91;94m \033[48;2;138;88;91m \033[48;2;138;86;90m \033[48;2;137;82;87m \033[48;2;139;80;86m \033[48;2;137;85;89m \033[48;2;137;85;89m \033[48;2;133;81;85m \033[48;2;143;90;95m \033[48;2;154;101;109m \033[48;2;163;110;122m \033[48;2;154;106;118m \033[48;2;160;112;123m \033[48;2;170;120;132m \033[48;2;165;118;130m \033[48;2;162;114;125m \033[48;2;158;110;122m \033[48;2;156;108;122m \033[48;2;156;108;122m \033[48;2;159;111;125m \033[48;2;156;112;122m \033[48;2;155;112;122m \033[48;2;153;110;120m \033[48;2;155;107;123m \033[48;2;153;96;117m \033[48;2;159;105;128m \033[48;2;181;138;161m \033[48;2;186;152;175m \033[48;2;178;154;177m \033[48;2;177;157;182m \033[48;2;177;157;182m \033[48;2;177;157;182m \033[48;2;180;160;185m \033[48;2;180;160;185m \033[48;2;177;158;182m \033[48;2;174;154;179m \033[48;2;171;151;176m \033[48;2;169;149;174m \033[48;2;166;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;164;151;180m \033[48;2;164;151;181m \033[48;2;163;150;180m \033[48;2;168;155;184m \033[48;2;171;158;188m \033[48;2;178;165;195m \033[48;2;178;165;195m \033[48;2;176;165;195m \033[48;2;176;165;195m \033[m");
$display("\033[48;2;176;165;197m \033[48;2;176;165;197m \033[48;2;177;163;196m \033[48;2;175;161;194m \033[48;2;175;161;194m \033[48;2;175;162;192m \033[48;2;179;166;196m \033[48;2;176;163;193m \033[48;2;173;158;189m \033[48;2;175;160;191m \033[48;2;175;160;191m \033[48;2;173;158;189m \033[48;2;171;156;187m \033[48;2;171;156;187m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;171;155;181m \033[48;2;171;155;181m \033[48;2;173;157;183m \033[48;2;183;163;188m \033[48;2;188;168;193m \033[48;2;186;166;192m \033[48;2;185;166;188m \033[48;2;186;167;189m \033[48;2;184;165;187m \033[48;2;177;158;177m \033[48;2;175;156;175m \033[48;2;179;160;179m \033[48;2;189;163;182m \033[48;2;188;160;180m \033[48;2;182;153;173m \033[48;2;185;145;158m \033[48;2;184;141;149m \033[48;2;160;107;113m \033[48;2;143;94;98m \033[48;2;143;94;98m \033[48;2;140;91;95m \033[48;2;140;90;93m \033[48;2;141;91;94m \033[48;2;138;88;91m \033[48;2;135;83;87m \033[48;2;134;80;85m \033[48;2;125;67;73m \033[48;2;121;61;67m \033[48;2;117;58;65m \033[48;2;115;58;63m \033[48;2;124;72;72m \033[48;2;121;69;72m \033[48;2;124;71;78m \033[48;2;125;72;80m \033[48;2;124;71;80m \033[48;2;142;89;97m \033[48;2;157;109;121m \033[48;2;160;113;125m \033[48;2;159;111;123m \033[48;2;158;111;120m \033[48;2;158;111;120m \033[48;2;159;112;121m \033[48;2;155;112;122m \033[48;2;155;112;122m \033[48;2;156;113;123m \033[48;2;161;114;130m \033[48;2;158;110;129m \033[48;2;181;144;162m \033[48;2;178;155;174m \033[48;2;181;160;179m \033[48;2;182;162;184m \033[48;2;182;162;187m \033[48;2;182;162;187m \033[48;2;176;156;181m \033[48;2;177;157;182m \033[48;2;182;162;187m \033[48;2;183;163;188m \033[48;2;183;163;188m \033[48;2;183;163;188m \033[48;2;175;155;180m \033[48;2;167;150;176m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;163;150;178m \033[48;2;163;150;180m \033[48;2;164;151;181m \033[48;2;173;160;190m \033[48;2;176;163;193m \033[48;2;178;165;195m \033[48;2;178;165;195m \033[48;2;177;166;196m \033[48;2;178;167;197m \033[m");
$display("\033[48;2;177;163;196m \033[48;2;176;162;195m \033[48;2;175;161;194m \033[48;2;175;161;194m \033[48;2;173;159;192m \033[48;2;173;159;192m \033[48;2;172;158;191m \033[48;2;172;158;191m \033[48;2;172;157;188m \033[48;2;172;157;188m \033[48;2;172;157;188m \033[48;2;171;156;187m \033[48;2;169;154;185m \033[48;2;170;155;186m \033[48;2;172;158;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;172;158;184m \033[48;2;172;158;184m \033[48;2;171;157;183m \033[48;2;175;155;183m \033[48;2;173;153;180m \033[48;2;179;159;184m \033[48;2;186;167;189m \033[48;2;187;168;190m \033[48;2;181;162;184m \033[48;2;182;163;185m \033[48;2;187;168;190m \033[48;2;186;167;189m \033[48;2;181;162;181m \033[48;2;181;162;181m \033[48;2;181;162;181m \033[48;2;185;164;183m \033[48;2;186;163;183m \033[48;2;183;158;179m \033[48;2;188;154;168m \033[48;2;177;136;146m \033[48;2;162;112;117m \033[48;2;141;91;90m \033[48;2;145;95;96m \033[48;2;142;91;96m \033[48;2;141;90;95m \033[48;2;141;91;94m \033[48;2;139;89;88m \033[48;2;137;87;90m \033[48;2;136;84;88m \033[48;2;137;80;86m \033[48;2;134;75;81m \033[48;2;129;70;76m \033[48;2;123;64;70m \033[48;2;118;68;72m \033[48;2;114;65;68m \033[48;2;103;54;57m \033[48;2;88;44;40m \033[48;2;87;41;40m \033[48;2;92;43;42m \033[48;2;114;59;65m \033[48;2;133;82;87m \033[48;2;154;103;113m \033[48;2;159;112;120m \033[48;2;159;112;120m \033[48;2;159;112;120m \033[48;2;155;113;115m \033[48;2;153;113;121m \033[48;2;152;115;128m \033[48;2;156;119;138m \033[48;2;187;154;173m \033[48;2;176;152;172m \033[48;2;173;153;176m \033[48;2;180;161;183m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;179;160;182m \033[48;2;175;155;180m \033[48;2;178;158;183m \033[48;2;182;162;187m \033[48;2;178;158;182m \033[48;2;177;158;180m \033[48;2;175;156;178m \033[48;2;170;150;176m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;167;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;152;176m \033[48;2;164;152;176m \033[48;2;163;151;175m \033[48;2;163;150;177m \033[48;2;163;150;180m \033[48;2;164;151;181m \033[48;2;166;153;183m \033[48;2;169;156;186m \033[48;2;170;157;187m \033[48;2;170;158;188m \033[48;2;172;161;191m \033[48;2;175;164;194m \033[m");
$display("\033[48;2;177;163;196m \033[48;2;177;163;196m \033[48;2;175;161;194m \033[48;2;175;161;194m \033[48;2;175;161;194m \033[48;2;174;161;191m \033[48;2;175;162;192m \033[48;2;175;162;192m \033[48;2;175;160;191m \033[48;2;174;159;190m \033[48;2;174;159;190m \033[48;2;171;157;183m \033[48;2;172;158;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;172;156;182m \033[48;2;172;156;182m \033[48;2;174;158;184m \033[48;2;183;163;188m \033[48;2;192;172;197m \033[48;2;193;173;198m \033[48;2;191;172;194m \033[48;2;190;171;193m \033[48;2;184;165;187m \033[48;2;188;169;191m \033[48;2;191;172;194m \033[48;2;191;172;194m \033[48;2;183;164;186m \033[48;2;185;166;186m \033[48;2;181;163;179m \033[48;2;189;168;187m \033[48;2;188;164;185m \033[48;2;187;162;183m \033[48;2;194;163;177m \033[48;2;170;127;136m \033[48;2;171;118;118m \033[48;2;157;108;103m \033[48;2;137;86;85m \033[48;2;142;92;95m \033[48;2;141;92;95m \033[48;2;142;93;96m \033[48;2;140;91;94m \033[48;2;141;91;94m \033[48;2;138;88;91m \033[48;2;135;85;88m \033[48;2;134;83;84m \033[48;2;134;77;83m \033[48;2;140;74;86m \033[48;2;147;82;95m \033[48;2;150;84;100m \033[48;2;146;77;99m \033[48;2;153;84;109m \033[48;2;156;93;113m \033[48;2;161;105;119m \033[48;2;162;112;124m \033[48;2;162;112;124m \033[48;2;158;108;120m \033[48;2;155;112;119m \033[48;2;155;112;119m \033[48;2;156;113;120m \033[48;2;152;118;119m \033[48;2;186;155;160m \033[48;2;184;161;170m \033[48;2;183;160;183m \033[48;2;183;159;183m \033[48;2;182;158;182m \033[48;2;178;156;179m \033[48;2;181;159;182m \033[48;2;184;162;185m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;179;160;182m \033[48;2;178;159;181m \033[48;2;178;159;181m \033[48;2;181;162;184m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;177;158;180m \033[48;2;172;153;175m \033[48;2;169;150;172m \033[48;2;168;148;173m \033[48;2;168;148;173m \033[48;2;169;149;174m \033[48;2;166;150;173m \033[48;2;165;150;173m \033[48;2;165;150;173m \033[48;2;165;149;174m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;170;157;183m \033[48;2;174;164;189m \033[48;2;178;168;193m \033[48;2;178;168;193m \033[48;2;177;167;192m \033[48;2;175;165;190m \033[m");
$display("\033[48;2;177;163;196m \033[48;2;177;163;196m \033[48;2;177;163;196m \033[48;2;177;163;196m \033[48;2;174;160;193m \033[48;2;173;160;190m \033[48;2;173;160;190m \033[48;2;173;160;190m \033[48;2;173;158;189m \033[48;2;173;158;189m \033[48;2;173;158;189m \033[48;2;171;157;183m \033[48;2;172;158;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;174;160;186m \033[48;2;174;160;186m \033[48;2;176;161;186m \033[48;2;176;160;187m \033[48;2;179;163;189m \033[48;2;186;166;191m \033[48;2;188;168;193m \033[48;2;190;170;195m \033[48;2;190;171;193m \033[48;2;188;169;191m \033[48;2;188;169;191m \033[48;2;185;166;188m \033[48;2;181;162;184m \033[48;2;184;165;187m \033[48;2;178;159;181m \033[48;2;182;163;182m \033[48;2;182;164;180m \033[48;2;186;165;184m \033[48;2;187;164;184m \033[48;2;182;156;178m \033[48;2;178;147;162m \033[48;2;170;125;134m \033[48;2;154;99;99m \033[48;2;160;111;107m \033[48;2;151;101;100m \033[48;2;143;93;96m \033[48;2;141;92;95m \033[48;2;141;92;95m \033[48;2;141;92;95m \033[48;2;141;91;94m \033[48;2;138;88;91m \033[48;2;136;86;89m \033[48;2;136;86;87m \033[48;2;134;77;83m \033[48;2;137;71;82m \033[48;2;133;68;82m \033[48;2;132;66;82m \033[48;2;140;74;93m \033[48;2;148;85;108m \033[48;2;155;99;116m \033[48;2;161;111;122m \033[48;2;157;114;124m \033[48;2;154;111;121m \033[48;2;155;112;122m \033[48;2;155;111;124m \033[48;2;155;111;124m \033[48;2;157;113;126m \033[48;2;182;150;164m \033[48;2;180;154;169m \033[48;2;180;159;179m \033[48;2;185;162;185m \033[48;2;185;161;185m \033[48;2;185;161;185m \033[48;2;181;159;183m \033[48;2;182;160;183m \033[48;2;180;158;181m \033[48;2;180;161;183m \033[48;2;180;161;183m \033[48;2;179;160;182m \033[48;2;177;158;180m \033[48;2;180;161;183m \033[48;2;181;162;184m \033[48;2;183;164;186m \033[48;2;183;164;186m \033[48;2;182;163;185m \033[48;2;179;160;182m \033[48;2;174;155;177m \033[48;2;172;153;175m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;166;150;173m \033[48;2;165;150;173m \033[48;2;165;150;173m \033[48;2;165;149;174m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;169;155;181m \033[48;2;174;161;187m \033[48;2;175;165;190m \033[48;2;177;167;192m \033[48;2;177;167;192m \033[48;2;176;166;191m \033[48;2;174;164;189m \033[m");
$display("\033[48;2;184;169;202m \033[48;2;176;161;194m \033[48;2;175;164;194m \033[48;2;172;161;191m \033[48;2;172;161;191m \033[48;2;174;160;185m \033[48;2;173;159;184m \033[48;2;173;159;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;182m \033[48;2;169;155;180m \033[48;2;172;158;183m \033[48;2;176;162;187m \033[48;2;175;161;186m \033[48;2;178;164;189m \033[48;2;185;165;190m \033[48;2;184;164;189m \033[48;2;185;165;190m \033[48;2;187;167;192m \033[48;2;187;167;192m \033[48;2;186;166;191m \033[48;2;183;164;186m \033[48;2;186;167;189m \033[48;2;186;167;189m \033[48;2;182;163;185m \033[48;2;182;163;185m \033[48;2;180;161;183m \033[48;2;176;157;175m \033[48;2;179;160;179m \033[48;2;178;159;178m \033[48;2;179;158;177m \033[48;2;180;157;177m \033[48;2;177;152;173m \033[48;2;180;145;167m \033[48;2;164;123;132m \033[48;2;148;99;99m \033[48;2;143;93;92m \033[48;2;144;94;93m \033[48;2;136;86;85m \033[48;2;136;87;90m \033[48;2;136;87;90m \033[48;2;136;87;90m \033[48;2;137;88;91m \033[48;2;137;88;91m \033[48;2;141;92;95m \033[48;2;139;93;94m \033[48;2;142;96;98m \033[48;2;151;103;109m \033[48;2;155;107;121m \033[48;2;158;110;126m \033[48;2;160;110;132m \033[48;2;163;111;132m \033[48;2;160;111;132m \033[48;2;157;112;131m \033[48;2;155;113;122m \033[48;2;152;110;120m \033[48;2;151;110;119m \033[48;2;154;108;123m \033[48;2;154;111;128m \033[48;2;157;121;138m \033[48;2;182;154;174m \033[48;2;179;156;176m \033[48;2;176;154;177m \033[48;2;177;155;178m \033[48;2;177;155;178m \033[48;2;176;154;177m \033[48;2;178;154;184m \033[48;2;178;155;183m \033[48;2;177;154;182m \033[48;2;175;155;180m \033[48;2;175;155;180m \033[48;2;175;155;180m \033[48;2;174;154;179m \033[48;2;179;159;184m \033[48;2;176;156;181m \033[48;2;174;156;177m \033[48;2;175;156;178m \033[48;2;176;157;179m \033[48;2;177;158;180m \033[48;2;174;155;177m \033[48;2;175;156;178m \033[48;2;176;156;181m \033[48;2;172;152;177m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;167;147;172m \033[48;2;169;149;174m \033[48;2;168;150;176m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;166;150;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;164;150;176m \033[48;2;165;151;177m \033[48;2;168;154;180m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;172;158;184m \033[48;2;173;158;185m \033[48;2;175;165;190m \033[48;2;177;167;192m \033[48;2;174;164;189m \033[48;2;174;164;189m \033[48;2;176;166;191m \033[m");
$display("\033[48;2;179;166;196m \033[48;2;176;163;193m \033[48;2;174;161;187m \033[48;2;173;160;186m \033[48;2;173;160;186m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;179;165;191m \033[48;2;174;160;185m \033[48;2;176;162;187m \033[48;2;174;160;185m \033[48;2;172;156;182m \033[48;2;174;158;184m \033[48;2;175;159;185m \033[48;2;178;158;183m \033[48;2;178;158;183m \033[48;2;178;158;183m \033[48;2;176;157;179m \033[48;2;174;155;177m \033[48;2;177;158;180m \033[48;2;178;159;181m \033[48;2;179;160;182m \033[48;2;178;159;181m \033[48;2;175;156;178m \033[48;2;176;157;179m \033[48;2;173;154;176m \033[48;2;175;154;173m \033[48;2;178;157;176m \033[48;2;176;155;174m \033[48;2;180;153;167m \033[48;2;168;130;142m \033[48;2;146;95;101m \033[48;2;144;91;95m \033[48;2;141;91;94m \033[48;2;135;86;89m \033[48;2;137;88;91m \033[48;2;136;87;90m \033[48;2;136;87;90m \033[48;2;137;87;90m \033[48;2;137;87;90m \033[48;2;136;86;89m \033[48;2;134;81;84m \033[48;2;136;84;90m \033[48;2;144;91;100m \033[48;2;152;97;106m \033[48;2;153;102;111m \033[48;2;156;105;117m \033[48;2;156;113;127m \033[48;2;157;112;129m \033[48;2;157;113;128m \033[48;2;153;109;124m \033[48;2;150;106;121m \033[48;2;151;107;122m \033[48;2;156;108;130m \033[48;2;153;110;130m \033[48;2;157;117;137m \033[48;2;187;154;177m \033[48;2;184;160;184m \033[48;2;184;159;185m \033[48;2;180;158;178m \033[48;2;180;159;178m \033[48;2;179;159;177m \033[48;2;176;153;179m \033[48;2;176;153;179m \033[48;2;178;155;181m \033[48;2;176;156;181m \033[48;2;176;156;181m \033[48;2;180;160;185m \033[48;2;180;160;185m \033[48;2;177;157;182m \033[48;2;176;156;181m \033[48;2;182;162;187m \033[48;2;182;162;187m \033[48;2;183;163;188m \033[48;2;182;162;187m \033[48;2;179;159;184m \033[48;2;175;155;180m \033[48;2;177;159;181m \033[48;2;180;161;183m \033[48;2;183;164;186m \033[48;2;181;161;187m \033[48;2;175;155;180m \033[48;2;169;149;174m \033[48;2;168;150;175m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;164;150;175m \033[48;2;164;150;175m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;177m \033[48;2;170;156;182m \033[48;2;177;163;189m \033[48;2;174;160;186m \033[48;2;177;164;190m \033[48;2;177;164;190m \033[48;2;175;162;188m \033[48;2;172;159;185m \033[48;2;171;158;184m \033[48;2;174;163;187m \033[48;2;177;167;192m \033[48;2;178;168;193m \033[m");
$display("\033[48;2;174;160;190m \033[48;2;174;160;190m \033[48;2;174;161;188m \033[48;2;173;161;187m \033[48;2;173;160;186m \033[48;2;173;159;184m \033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;171;157;183m \033[48;2;172;158;184m \033[48;2;171;157;183m \033[48;2;168;154;180m \033[48;2;166;152;178m \033[48;2;168;154;180m \033[48;2;166;152;177m \033[48;2;166;152;177m \033[48;2;166;152;177m \033[48;2;166;151;176m \033[48;2;166;151;176m \033[48;2;166;151;176m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;168;148;173m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;169;150;172m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;146;167m \033[48;2;169;149;167m \033[48;2;167;147;165m \033[48;2;173;144;160m \033[48;2;171;134;146m \033[48;2;146;94;99m \033[48;2;141;87;93m \033[48;2;137;86;90m \033[48;2;140;91;94m \033[48;2;137;88;91m \033[48;2;137;88;91m \033[48;2;137;88;91m \033[48;2;137;87;90m \033[48;2;136;86;89m \033[48;2;133;83;86m \033[48;2;131;80;76m \033[48;2;128;77;74m \033[48;2;130;78;80m \033[48;2;131;78;80m \033[48;2;130;81;84m \033[48;2;140;90;94m \033[48;2;136;94;102m \033[48;2;139;96;105m \033[48;2;143;100;110m \033[48;2;146;102;118m \033[48;2;155;111;126m \033[48;2;154;109;125m \033[48;2;159;106;129m \033[48;2;154;104;126m \033[48;2;140;95;116m \033[48;2;101;66;77m \033[48;2;138;110;122m \033[48;2;182;154;169m \033[48;2;175;153;171m \033[48;2;175;154;172m \033[48;2;174;153;172m \033[48;2;172;150;174m \033[48;2;172;150;175m \033[48;2;172;149;175m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;170;151;175m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;170;150;175m \033[48;2;170;149;175m \033[48;2;171;149;175m \033[48;2;169;149;173m \033[48;2;172;152;177m \033[48;2;172;152;177m \033[48;2;170;151;175m \033[48;2;171;152;174m \033[48;2;171;152;174m \033[48;2;170;151;173m \033[48;2;168;149;173m \033[48;2;168;150;174m \033[48;2;169;150;174m \033[48;2;166;150;175m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;162;149;174m \033[48;2;165;151;177m \033[48;2;163;150;176m \033[48;2;164;151;177m \033[48;2;162;149;175m \033[48;2;162;149;175m \033[48;2;163;151;177m \033[48;2;161;151;176m \033[48;2;162;153;179m \033[m");
$display("\033[48;2;171;156;187m \033[48;2;171;156;187m \033[48;2;170;155;186m \033[48;2;171;156;187m \033[48;2;171;156;187m \033[48;2;170;155;186m \033[48;2;170;155;186m \033[48;2;170;155;186m \033[48;2;170;156;182m \033[48;2;169;155;181m \033[48;2;166;152;178m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;166;151;174m \033[48;2;166;151;174m \033[48;2;166;151;174m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;168;148;173m \033[48;2;167;148;170m \033[48;2;167;148;170m \033[48;2;167;148;170m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;169;150;172m \033[48;2;170;149;168m \033[48;2;172;148;165m \033[48;2;174;147;162m \033[48;2;177;147;148m \033[48;2;174;133;136m \033[48;2;147;90;98m \033[48;2;146;87;93m \033[48;2;141;85;91m \033[48;2;138;86;90m \033[48;2;137;88;91m \033[48;2;137;88;91m \033[48;2;137;88;91m \033[48;2;137;87;90m \033[48;2;134;84;87m \033[48;2;133;83;86m \033[48;2;128;78;81m \033[48;2;127;78;80m \033[48;2;132;82;85m \033[48;2;137;86;91m \033[48;2;139;88;97m \033[48;2;150;99;111m \033[48;2;149;101;115m \033[48;2;151;102;121m \033[48;2;155;106;127m \033[48;2;159;104;129m \033[48;2;159;106;129m \033[48;2;161;105;130m \033[48;2;162;108;129m \033[48;2;158;111;131m \033[48;2;173;137;155m \033[48;2;134;102;123m \033[48;2;87;58;74m \033[48;2;84;61;72m \033[48;2;102;85;86m \033[48;2;149;129;131m \033[48;2;181;162;165m \033[48;2;175;155;170m \033[48;2;176;155;173m \033[48;2;175;154;173m \033[48;2;175;153;176m \033[48;2;175;153;176m \033[48;2;175;153;176m \033[48;2;169;151;176m \033[48;2;171;151;176m \033[48;2;171;151;176m \033[48;2;170;151;173m \033[48;2;170;151;173m \033[48;2;169;150;172m \033[48;2;170;151;173m \033[48;2;170;151;173m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;168;151;177m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;167;151;177m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;166;152;177m \033[48;2;164;150;175m \033[48;2;163;151;175m \033[48;2;163;151;175m \033[48;2;163;150;177m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[48;2;162;150;178m \033[48;2;160;149;179m \033[48;2;160;149;179m \033[m");
$display("\033[48;2;173;159;185m \033[48;2;173;159;185m \033[48;2;172;158;184m \033[48;2;171;157;183m \033[48;2;171;157;183m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;170;156;182m \033[48;2;169;155;181m \033[48;2;169;155;181m \033[48;2;166;152;175m \033[48;2;170;156;179m \033[48;2;171;157;180m \033[48;2;176;161;182m \033[48;2;178;163;184m \033[48;2;175;160;181m \033[48;2;176;157;179m \033[48;2;176;157;179m \033[48;2;178;159;181m \033[48;2;178;159;181m \033[48;2;178;159;181m \033[48;2;177;158;180m \033[48;2;173;154;173m \033[48;2;173;154;173m \033[48;2;174;155;174m \033[48;2;176;157;176m \033[48;2;175;156;175m \033[48;2;175;156;175m \033[48;2;170;156;173m \033[48;2;175;158;175m \033[48;2;173;153;171m \033[48;2;171;149;166m \033[48;2;181;152;165m \033[48;2;184;147;158m \033[48;2;176;130;130m \033[48;2;204;153;153m \033[48;2;164;114;116m \033[48;2;154;109;113m \033[48;2;149;105;108m \033[48;2;145;104;108m \033[48;2;144;105;108m \033[48;2;139;101;103m \033[48;2;137;98;99m \033[48;2;132;90;94m \033[48;2;127;82;86m \033[48;2;133;82;87m \033[48;2;147;96;100m \033[48;2;148;97;104m \033[48;2;151;100;108m \033[48;2;156;102;116m \033[48;2;159;105;123m \033[48;2;159;103;125m \033[48;2;160;102;127m \033[48;2;160;102;127m \033[48;2;160;102;127m \033[48;2;161;101;127m \033[48;2;161;101;127m \033[48;2;162;102;128m \033[48;2;157;103;127m \033[48;2;149;107;126m \033[48;2;167;136;156m \033[48;2;152;131;156m \033[48;2;80;61;84m \033[48;2;79;60;80m \033[48;2;70;56;65m \033[48;2;73;61;64m \033[48;2;79;68;66m \033[48;2;112;96;93m \033[48;2;144;125;126m \033[48;2;161;135;148m \033[48;2;173;152;163m \033[48;2;179;157;170m \033[48;2;177;155;170m \033[48;2;176;155;170m \033[48;2;176;155;172m \033[48;2;175;153;174m \033[48;2;172;153;172m \033[48;2;171;154;172m \033[48;2;170;153;171m \033[48;2;171;152;171m \033[48;2;171;152;171m \033[48;2;170;151;170m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;170;151;173m \033[48;2;168;150;174m \033[48;2;166;151;174m \033[48;2;166;151;174m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;176m \033[48;2;165;151;177m \033[48;2;167;153;179m \033[48;2;173;159;185m \033[48;2;173;159;184m \033[48;2;175;161;186m \033[48;2;177;163;188m \033[48;2;178;164;189m \033[48;2;178;164;189m \033[48;2;178;164;189m \033[48;2;176;164;188m \033[48;2;174;162;186m \033[48;2;173;161;185m \033[m");
$display("\033[48;2;175;161;187m \033[48;2;175;161;187m \033[48;2;173;159;185m \033[48;2;172;158;184m \033[48;2;170;156;182m \033[48;2;168;153;179m \033[48;2;166;150;176m \033[48;2;168;152;178m \033[48;2;168;153;179m \033[48;2;166;152;178m \033[48;2;166;151;177m \033[48;2;165;150;174m \033[48;2;175;160;182m \033[48;2;178;164;184m \033[48;2;183;168;187m \033[48;2;183;166;185m \033[48;2;180;163;183m \033[48;2;182;163;183m \033[48;2;186;167;186m \033[48;2;185;166;185m \033[48;2;184;166;184m \033[48;2;186;166;186m \033[48;2;186;167;187m \033[48;2;179;163;180m \033[48;2;177;160;177m \033[48;2;183;163;182m \033[48;2;183;165;183m \033[48;2;181;164;181m \033[48;2;175;158;174m \033[48;2;172;151;166m \033[48;2;171;148;159m \033[48;2;165;138;144m \033[48;2;177;146;151m \033[48;2;195;159;164m \033[48;2;173;128;133m \033[48;2;172;130;133m \033[48;2;119;83;85m \033[48;2;143;112;111m \033[48;2;143;124;133m \033[48;2;133;115;123m \033[48;2;149;137;145m \033[48;2;146;128;139m \033[48;2;150;133;146m \033[48;2;135;117;132m \033[48;2;147;127;140m \033[48;2;144;115;125m \033[48;2;128;88;96m \033[48;2;136;83;92m \033[48;2;144;91;99m \033[48;2;147;96;104m \033[48;2;151;96;109m \033[48;2;152;95;114m \033[48;2;154;96;118m \033[48;2;159;97;121m \033[48;2;161;98;123m \033[48;2;162;99;126m \033[48;2;162;100;126m \033[48;2;160;100;126m \033[48;2;158;100;125m \033[48;2;141;91;112m \033[48;2;163;126;145m \033[48;2;168;144;166m \033[48;2;154;138;161m \033[48;2;80;62;85m \033[48;2;77;60;79m \033[48;2;68;55;65m \033[48;2;68;56;60m \033[48;2;65;55;54m \033[48;2;64;54;52m \033[48;2;74;58;58m \033[48;2;105;85;81m \033[48;2;120;90;90m \033[48;2;130;99;101m \033[48;2;136;102;107m \033[48;2;138;108;112m \033[48;2;135;105;112m \033[48;2;147;118;125m \033[48;2;155;129;140m \033[48;2;169;142;151m \033[48;2;177;150;160m \033[48;2;180;160;174m \033[48;2;179;160;177m \033[48;2;177;156;178m \033[48;2;177;156;177m \033[48;2;175;155;175m \033[48;2;176;159;178m \033[48;2;176;159;178m \033[48;2;176;159;179m \033[48;2;177;158;180m \033[48;2;173;156;176m \033[48;2;171;155;174m \033[48;2;168;151;175m \033[48;2;167;151;175m \033[48;2;167;151;175m \033[48;2;167;151;175m \033[48;2;166;151;177m \033[48;2;166;151;177m \033[48;2;166;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;152;178m \033[48;2;169;155;181m \033[48;2;172;158;184m \033[48;2;177;163;188m \033[48;2;178;165;190m \033[48;2;177;165;189m \033[48;2;176;163;188m \033[48;2;175;163;187m \033[48;2;173;161;185m \033[48;2;174;162;186m \033[m");
$display("\033[48;2;174;160;186m \033[48;2;174;160;186m \033[48;2;171;157;183m \033[48;2;170;156;182m \033[48;2;167;153;179m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;165;149;175m \033[48;2;166;150;176m \033[48;2;172;157;179m \033[48;2;176;161;179m \033[48;2;179;160;179m \033[48;2;181;162;181m \033[48;2;178;159;178m \033[48;2;177;158;177m \033[48;2;182;163;182m \033[48;2;180;161;180m \033[48;2;180;162;178m \033[48;2;182;164;180m \033[48;2;179;161;177m \033[48;2;174;157;169m \033[48;2;171;151;163m \033[48;2;164;140;154m \033[48;2;161;128;140m \033[48;2;157;124;133m \033[48;2;162;129;135m \033[48;2;160;129;130m \033[48;2;164;128;128m \033[48;2;161;125;124m \033[48;2;193;158;162m \033[48;2;167;132;137m \033[48;2;167;126;132m \033[48;2;147;106;110m \033[48;2;139;103;105m \033[48;2;121;91;91m \033[48;2;122;104;102m \033[48;2;114;99;99m \033[48;2;114;102;105m \033[48;2;123;106;112m \033[48;2;112;95;104m \033[48;2;113;95;110m \033[48;2;121;101;113m \033[48;2;120;92;101m \033[48;2;125;82;91m \033[48;2;128;75;83m \033[48;2;131;78;86m \033[48;2;138;85;93m \033[48;2;144;87;96m \033[48;2;147;89;101m \033[48;2;151;93;108m \033[48;2;155;94;109m \033[48;2;158;97;115m \033[48;2;162;100;122m \033[48;2;161;98;117m \033[48;2;147;92;108m \033[48;2;135;90;103m \033[48;2;158;130;143m \033[48;2;163;145;159m \033[48;2;166;148;170m \033[48;2;149;128;154m \033[48;2;79;60;82m \033[48;2;75;56;76m \033[48;2;66;53;62m \033[48;2;65;54;58m \033[48;2;64;54;55m \033[48;2;58;52;50m \033[48;2;61;51;49m \033[48;2;63;51;43m \033[48;2;84;61;56m \033[48;2;111;85;80m \033[48;2;115;84;82m \033[48;2;112;81;80m \033[48;2;108;77;76m \033[48;2;113;82;81m \033[48;2;116;85;81m \033[48;2;125;93;90m \033[48;2;131;100;97m \033[48;2;135;107;104m \033[48;2;132;105;102m \033[48;2;135;105;107m \033[48;2;140;106;118m \033[48;2;146;116;127m \033[48;2;152;125;135m \033[48;2;163;140;148m \033[48;2;174;153;161m \033[48;2;178;154;167m \033[48;2;179;160;177m \033[48;2;174;156;173m \033[48;2;172;153;172m \033[48;2;169;151;174m \033[48;2;167;152;175m \033[48;2;167;152;175m \033[48;2;167;151;177m \033[48;2;167;151;177m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;166;152;178m \033[48;2;168;156;180m \033[48;2;172;160;184m \033[48;2;172;160;184m \033[48;2;172;160;184m \033[48;2;172;160;184m \033[48;2;173;161;185m \033[m");
$display("\033[48;2;171;155;182m \033[48;2;171;155;182m \033[48;2;170;154;180m \033[48;2;170;154;180m \033[48;2;167;151;177m \033[48;2;168;152;178m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;151;174m \033[48;2;165;150;173m \033[48;2;165;150;173m \033[48;2;168;153;174m \033[48;2;173;158;179m \033[48;2;176;161;182m \033[48;2;181;162;181m \033[48;2;185;166;185m \033[48;2;180;161;180m \033[48;2;176;160;179m \033[48;2;182;164;181m \033[48;2;175;153;168m \033[48;2;172;147;164m \033[48;2;164;136;148m \033[48;2;160;129;136m \033[48;2;153;124;127m \033[48;2;145;113;116m \033[48;2;140;105;104m \033[48;2;134;95;100m \033[48;2;135;99;100m \033[48;2;130;99;98m \033[48;2;142;111;106m \033[48;2;145;114;109m \033[48;2;170;139;134m \033[48;2;188;153;154m \033[48;2;164;129;135m \033[48;2;158;122;134m \033[48;2;131;96;102m \033[48;2;129;98;99m \033[48;2;123;96;88m \033[48;2;116;98;94m \033[48;2;117;102;100m \033[48;2;115;103;104m \033[48;2;118;101;109m \033[48;2;125;108;116m \033[48;2;122;105;113m \033[48;2;128;113;122m \033[48;2;126;97;108m \033[48;2;126;80;93m \033[48;2;131;73;85m \033[48;2;131;73;85m \033[48;2;135;77;89m \033[48;2;140;83;91m \033[48;2;143;86;95m \033[48;2;147;90;99m \033[48;2;151;90;107m \033[48;2;155;94;110m \033[48;2;144;83;99m \033[48;2;127;75;88m \033[48;2;140;96;114m \033[48;2;161;129;150m \033[48;2;167;145;172m \033[48;2;161;145;174m \033[48;2;166;148;175m \033[48;2;138;119;142m \033[48;2;79;60;78m \033[48;2;75;58;69m \033[48;2;66;56;58m \033[48;2;64;54;53m \033[48;2;62;52;49m \033[48;2;58;51;45m \033[48;2;58;51;43m \033[48;2;55;48;38m \033[48;2;59;46;36m \033[48;2;60;46;38m \033[48;2;78;60;53m \033[48;2;97;75;70m \033[48;2;92;68;64m \033[48;2;99;70;68m \033[48;2;99;69;67m \033[48;2;105;75;73m \033[48;2;109;79;77m \033[48;2;108;78;76m \033[48;2;105;75;73m \033[48;2;108;78;76m \033[48;2;110;79;80m \033[48;2;114;83;83m \033[48;2;112;81;81m \033[48;2;110;80;80m \033[48;2;113;83;83m \033[48;2;115;85;85m \033[48;2;122;94;94m \033[48;2;126;96;99m \033[48;2;134;109;113m \033[48;2;153;130;142m \033[48;2;170;146;163m \033[48;2;173;155;174m \033[48;2;171;154;173m \033[48;2;171;153;175m \033[48;2;169;151;177m \033[48;2;168;151;174m \033[48;2;166;151;173m \033[48;2;166;150;177m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;151;177m \033[48;2;164;151;177m \033[48;2;163;150;176m \033[48;2;161;150;175m \033[48;2;164;154;179m \033[48;2;167;157;182m \033[m");
$display("\033[48;2;171;155;182m \033[48;2;168;152;179m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;168;149;171m \033[48;2;168;149;172m \033[48;2;168;149;172m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;170;149;172m \033[48;2;172;153;175m \033[48;2;173;154;177m \033[48;2;178;157;177m \033[48;2;174;152;168m \033[48;2;167;143;157m \033[48;2;159;139;143m \033[48;2;160;132;135m \033[48;2;159;124;126m \033[48;2;151;112;117m \033[48;2;132;92;94m \033[48;2;124;86;85m \033[48;2;122;87;78m \033[48;2;100;66;56m \033[48;2;95;62;53m \033[48;2;100;72;63m \033[48;2;91;64;53m \033[48;2;100;75;62m \033[48;2;121;100;81m \033[48;2;136;113;97m \033[48;2;180;152;141m \033[48;2;175;146;142m \033[48;2;158;133;136m \033[48;2;152;131;139m \033[48;2;131;105;114m \033[48;2;142;114;119m \033[48;2;120;89;89m \033[48;2;118;100;98m \033[48;2;115;100;101m \033[48;2;112;102;103m \033[48;2;114;102;108m \033[48;2;113;101;108m \033[48;2;117;103;110m \033[48;2;128;111;120m \033[48;2;131;98;111m \033[48;2;132;83;102m \033[48;2;135;77;92m \033[48;2;135;77;92m \033[48;2;134;76;91m \033[48;2;138;81;90m \033[48;2;142;85;94m \033[48;2;141;84;93m \033[48;2;141;79;85m \033[48;2;129;73;85m \033[48;2;138;90;111m \033[48;2;154;128;144m \033[48;2;156;135;156m \033[48;2;160;145;174m \033[48;2;163;148;177m \033[48;2;164;148;175m \033[48;2;169;150;175m \033[48;2;129;110;129m \033[48;2;74;55;70m \033[48;2;70;53;61m \033[48;2;64;55;54m \033[48;2;61;53;50m \033[48;2;59;52;44m \033[48;2;57;50;40m \033[48;2;57;51;39m \033[48;2;57;51;36m \033[48;2;53;48;28m \033[48;2;53;48;29m \033[48;2;52;47;28m \033[48;2;59;48;34m \033[48;2;75;59;47m \033[48;2;84;65;54m \033[48;2;88;66;60m \033[48;2;89;65;59m \033[48;2;86;63;56m \033[48;2;81;57;53m \033[48;2;83;60;55m \033[48;2;84;60;55m \033[48;2;83;60;57m \033[48;2;83;60;57m \033[48;2;80;56;53m \033[48;2;82;57;56m \033[48;2;88;63;61m \033[48;2;84;61;59m \033[48;2;90;66;65m \033[48;2;99;76;74m \033[48;2;106;82;80m \033[48;2;113;85;87m \033[48;2;120;90;92m \033[48;2;122;92;95m \033[48;2;114;87;90m \033[48;2;125;98;102m \033[48;2;132;112;115m \033[48;2;158;138;143m \033[48;2;171;155;165m \033[48;2;170;154;171m \033[48;2;166;151;171m \033[48;2;166;151;173m \033[48;2;166;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[m");
$display("\033[48;2;171;155;182m \033[48;2;171;155;182m \033[48;2;169;153;179m \033[48;2;169;153;179m \033[48;2;165;149;175m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;167;148;170m \033[48;2;167;148;170m \033[48;2;167;148;170m \033[48;2;167;149;166m \033[48;2;169;144;163m \033[48;2;168;138;158m \033[48;2;159;130;140m \033[48;2;162;130;138m \033[48;2;155;121;128m \033[48;2;144;109;112m \033[48;2;128;93;92m \033[48;2;108;74;70m \033[48;2;96;65;64m \033[48;2;85;54;47m \033[48;2;79;48;37m \033[48;2;66;45;32m \033[48;2;83;62;48m \033[48;2;84;62;49m \033[48;2;71;51;40m \033[48;2;71;52;38m \033[48;2;76;56;42m \033[48;2;114;92;73m \033[48;2;135;112;96m \033[48;2;185;157;146m \033[48;2;171;141;143m \033[48;2;163;136;145m \033[48;2;165;142;160m \033[48;2;133;113;121m \033[48;2;125;102;106m \033[48;2;120;93;93m \033[48;2;115;97;95m \033[48;2;112;97;97m \033[48;2;118;106;108m \033[48;2;117;104;110m \033[48;2;117;104;110m \033[48;2;116;103;110m \033[48;2;133;115;123m \033[48;2;138;106;120m \033[48;2;129;80;99m \033[48;2;129;71;86m \033[48;2;129;71;86m \033[48;2;130;72;87m \033[48;2;129;72;81m \033[48;2;130;73;82m \033[48;2;130;73;82m \033[48;2;134;89;101m \033[48;2;157;123;140m \033[48;2;153;136;157m \033[48;2;156;143;173m \033[48;2;158;145;173m \033[48;2;162;148;177m \033[48;2;164;149;178m \033[48;2;162;145;171m \033[48;2;164;145;170m \033[48;2;86;68;88m \033[48;2;73;55;67m \033[48;2;67;50;57m \033[48;2;61;53;51m \033[48;2;58;50;48m \033[48;2;58;51;43m \033[48;2;57;50;40m \033[48;2;57;51;39m \033[48;2;57;51;36m \033[48;2;54;49;29m \033[48;2;51;46;27m \033[48;2;50;45;26m \033[48;2;50;44;28m \033[48;2;54;46;30m \033[48;2;62;50;37m \033[48;2;76;58;51m \033[48;2;78;62;53m \033[48;2;76;60;52m \033[48;2;75;58;51m \033[48;2;75;58;51m \033[48;2;73;56;48m \033[48;2;68;51;47m \033[48;2;69;51;47m \033[48;2;69;51;47m \033[48;2;67;49;45m \033[48;2;68;50;46m \033[48;2;69;51;47m \033[48;2;69;51;47m \033[48;2;69;51;47m \033[48;2;73;54;51m \033[48;2;74;58;56m \033[48;2;68;51;50m \033[48;2;67;51;48m \033[48;2;74;53;55m \033[48;2;70;50;52m \033[48;2;68;52;51m \033[48;2;72;54;56m \033[48;2;77;59;70m \033[48;2;120;102;120m \033[48;2;170;156;175m \033[48;2;169;154;175m \033[48;2;166;150;176m \033[48;2;165;151;177m \033[48;2;165;151;177m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[48;2;163;150;176m \033[48;2;163;150;176m \033[m");
$display("\033[48;2;171;156;179m \033[48;2;170;155;178m \033[48;2;171;151;176m \033[48;2;169;149;174m \033[48;2;169;149;174m \033[48;2;168;149;170m \033[48;2;166;149;168m \033[48;2;169;151;166m \033[48;2;165;144;162m \033[48;2;163;139;155m \033[48;2;161;133;149m \033[48;2;155;123;138m \033[48;2;151;114;128m \033[48;2;146;108;118m \033[48;2;138;96;105m \033[48;2;124;85;89m \033[48;2;110;70;71m \033[48;2;91;56;54m \033[48;2;76;50;41m \033[48;2;66;48;34m \033[48;2;65;49;34m \033[48;2;62;49;33m \033[48;2;60;50;34m \033[48;2;63;51;36m \033[48;2;60;48;32m \033[48;2;63;51;35m \033[48;2;62;51;35m \033[48;2;63;51;35m \033[48;2;67;55;40m \033[48;2;96;80;62m \033[48;2;127;106;87m \033[48;2;185;158;150m \033[48;2;171;141;141m \033[48;2;154;129;137m \033[48;2;158;136;153m \033[48;2;126;103;117m \033[48;2;122;101;106m \033[48;2;115;96;92m \033[48;2;112;97;91m \033[48;2;115;99;99m \033[48;2;116;101;106m \033[48;2;114;101;111m \033[48;2;116;103;111m \033[48;2;111;99;103m \033[48;2;133;114;122m \033[48;2;139;106;119m \033[48;2;125;76;95m \033[48;2;129;66;83m \033[48;2;131;67;84m \033[48;2;126;69;84m \033[48;2;125;72;86m \033[48;2;135;92;107m \033[48;2;156;126;144m \033[48;2;153;131;151m \033[48;2;155;140;163m \033[48;2;158;149;176m \033[48;2;162;147;178m \033[48;2;162;147;178m \033[48;2;162;147;178m \033[48;2;161;145;172m \033[48;2;161;144;168m \033[48;2;94;75;90m \033[48;2;74;58;66m \033[48;2;68;53;57m \033[48;2;62;52;51m \033[48;2;60;50;48m \033[48;2;60;51;44m \033[48;2;60;51;42m \033[48;2;55;53;35m \033[48;2;54;51;34m \033[48;2;53;50;33m \033[48;2;53;50;31m \033[48;2;52;49;30m \033[48;2;50;47;28m \033[48;2;48;46;27m \033[48;2;49;44;25m \033[48;2;53;44;27m \033[48;2;55;42;26m \033[48;2;66;53;38m \033[48;2;71;57;46m \033[48;2;75;61;52m \033[48;2;72;58;49m \033[48;2;70;56;47m \033[48;2;65;54;45m \033[48;2;63;53;44m \033[48;2;60;50;41m \033[48;2;58;49;42m \033[48;2;58;49;42m \033[48;2;56;47;41m \033[48;2;55;47;40m \033[48;2;54;48;40m \033[48;2;56;49;42m \033[48;2;56;50;45m \033[48;2;53;48;46m \033[48;2;59;54;56m \033[48;2;58;54;57m \033[48;2;61;56;60m \033[48;2;64;59;63m \033[48;2;65;59;67m \033[48;2;70;62;72m \033[48;2;74;63;75m \033[48;2;106;90;106m \033[48;2;169;154;173m \033[48;2;168;153;174m \033[48;2;166;151;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;164;150;176m \033[48;2;164;150;176m \033[m");
$display("\033[48;2;172;157;180m \033[48;2;169;154;177m \033[48;2;166;151;172m \033[48;2;168;149;171m \033[48;2;170;148;171m \033[48;2;174;146;173m \033[48;2;150;122;138m \033[48;2;152;121;130m \033[48;2;145;113;119m \033[48;2;142;109;115m \033[48;2;130;99;104m \033[48;2;127;87;89m \033[48;2;117;82;82m \033[48;2;100;69;67m \033[48;2;85;57;47m \033[48;2;76;52;42m \033[48;2;67;46;35m \033[48;2;60;51;36m \033[48;2;60;51;36m \033[48;2;59;50;35m \033[48;2;58;51;33m \033[48;2;58;51;30m \033[48;2;58;52;28m \033[48;2;58;51;32m \033[48;2;58;51;32m \033[48;2;59;52;33m \033[48;2;62;55;37m \033[48;2;63;56;38m \033[48;2;64;57;39m \033[48;2;82;66;47m \033[48;2;131;107;88m \033[48;2;187;158;150m \033[48;2;168;138;138m \033[48;2;152;126;133m \033[48;2;151;128;144m \033[48;2;113;93;99m \033[48;2;108;88;90m \033[48;2;113;93;88m \033[48;2;109;98;94m \033[48;2;112;101;99m \033[48;2;113;101;103m \033[48;2;113;100;107m \033[48;2;116;103;110m \033[48;2;115;102;109m \033[48;2;123;109;113m \033[48;2;138;107;118m \033[48;2;121;73;89m \033[48;2;127;70;81m \033[48;2;127;84;96m \033[48;2;136;107;122m \033[48;2;144;128;146m \033[48;2;141;130;147m \033[48;2;151;139;160m \033[48;2;152;142;167m \033[48;2;155;145;170m \033[48;2;158;148;173m \033[48;2;160;148;179m \033[48;2;159;144;173m \033[48;2;158;142;168m \033[48;2;150;134;161m \033[48;2;78;65;76m \033[48;2;69;57;56m \033[48;2;63;56;50m \033[48;2;63;56;50m \033[48;2;59;52;46m \033[48;2;59;52;44m \033[48;2;59;52;42m \033[48;2;58;52;39m \033[48;2;53;50;33m \033[48;2;53;50;33m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;50;47;30m \033[48;2;51;50;30m \033[48;2;49;46;27m \033[48;2;50;43;25m \033[48;2;55;46;32m \033[48;2;56;46;31m \033[48;2;68;58;44m \033[48;2;92;77;68m \033[48;2;77;62;53m \033[48;2;67;53;44m \033[48;2;56;49;39m \033[48;2;56;49;39m \033[48;2;55;48;38m \033[48;2;54;51;38m \033[48;2;54;50;37m \033[48;2;55;51;41m \033[48;2;59;51;48m \033[48;2;59;51;48m \033[48;2;59;51;48m \033[48;2;57;53;52m \033[48;2;55;53;54m \033[48;2;59;57;58m \033[48;2;62;60;62m \033[48;2;62;60;63m \033[48;2;63;61;64m \033[48;2;64;61;66m \033[48;2;62;59;68m \033[48;2;64;60;75m \033[48;2;72;66;81m \033[48;2;115;104;122m \033[48;2;170;154;176m \033[48;2;168;151;176m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;149;176m \033[48;2;165;149;176m \033[m");
$display("\033[48;2;170;155;178m \033[48;2;167;152;175m \033[48;2;166;151;172m \033[48;2;168;149;171m \033[48;2;170;148;171m \033[48;2;130;97;119m \033[48;2;121;88;101m \033[48;2;116;80;85m \033[48;2;104;73;74m \033[48;2;96;63;65m \033[48;2;88;56;57m \033[48;2;81;55;51m \033[48;2;72;51;47m \033[48;2;70;53;45m \033[48;2;68;53;40m \033[48;2;62;52;37m \033[48;2;60;53;37m \033[48;2;60;51;36m \033[48;2;60;51;36m \033[48;2;60;51;36m \033[48;2;58;51;33m \033[48;2;58;51;30m \033[48;2;58;52;28m \033[48;2;58;51;32m \033[48;2;58;51;32m \033[48;2;60;53;34m \033[48;2;61;54;36m \033[48;2;61;54;36m \033[48;2;64;57;39m \033[48;2;78;61;43m \033[48;2;137;115;97m \033[48;2;182;153;145m \033[48;2;159;128;133m \033[48;2;149;121;136m \033[48;2;146;122;144m \033[48;2;110;87;102m \033[48;2;102;82;91m \033[48;2;117;97;99m \033[48;2;116;104;105m \033[48;2;113;102;106m \033[48;2;106;93;102m \033[48;2;115;102;109m \033[48;2;105;92;99m \033[48;2;114;102;108m \033[48;2;120;107;117m \033[48;2;147;127;138m \033[48;2;142;113;128m \033[48;2;145;125;137m \033[48;2;144;127;143m \033[48;2;147;133;153m \033[48;2;152;133;156m \033[48;2;152;138;163m \033[48;2;156;143;171m \033[48;2;154;144;169m \033[48;2;157;147;172m \033[48;2;156;146;171m \033[48;2;157;146;176m \033[48;2;157;142;172m \033[48;2;134;118;144m \033[48;2;78;66;76m \033[48;2;66;54;59m \033[48;2;63;52;50m \033[48;2;62;55;49m \033[48;2;62;55;49m \033[48;2;59;52;46m \033[48;2;59;52;44m \033[48;2;59;52;42m \033[48;2;57;51;38m \033[48;2;53;50;33m \033[48;2;53;50;33m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;51;50;30m \033[48;2;52;49;30m \033[48;2;54;47;29m \033[48;2;52;46;31m \033[48;2;54;49;33m \033[48;2;52;47;32m \033[48;2;53;45;34m \033[48;2;56;48;37m \033[48;2;55;45;35m \033[48;2;54;47;37m \033[48;2;52;45;35m \033[48;2;55;48;38m \033[48;2;54;50;41m \033[48;2;57;52;45m \033[48;2;59;54;50m \033[48;2;62;58;59m \033[48;2;60;58;59m \033[48;2;59;57;58m \033[48;2;56;53;55m \033[48;2;56;55;56m \033[48;2;62;60;61m \033[48;2;62;59;62m \033[48;2;62;60;63m \033[48;2;63;61;64m \033[48;2;63;60;65m \033[48;2;63;60;69m \033[48;2;64;60;75m \033[48;2;68;61;76m \033[48;2;85;74;91m \033[48;2;159;144;165m \033[48;2;168;151;177m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;149;176m \033[48;2;164;148;175m \033[m");
$display("\033[48;2;167;152;173m \033[48;2;166;151;172m \033[48;2;168;149;171m \033[48;2;169;151;173m \033[48;2;158;131;156m \033[48;2;88;57;72m \033[48;2;83;55;59m \033[48;2;77;49;43m \033[48;2;75;51;45m \033[48;2;73;54;45m \033[48;2;63;53;42m \033[48;2;62;53;38m \033[48;2;60;51;36m \033[48;2;69;60;45m \033[48;2;69;60;43m \033[48;2;61;52;35m \033[48;2;61;52;35m \033[48;2;60;51;34m \033[48;2;58;49;32m \033[48;2;58;49;32m \033[48;2;56;49;31m \033[48;2;56;49;31m \033[48;2;56;49;31m \033[48;2;56;51;31m \033[48;2;57;52;32m \033[48;2;58;53;33m \033[48;2;59;52;33m \033[48;2;62;55;36m \033[48;2;64;57;38m \033[48;2;72;62;37m \033[48;2;125;108;86m \033[48;2;159;134;126m \033[48;2;148;120;129m \033[48;2;150;125;138m \033[48;2;147;124;141m \033[48;2;162;142;154m \033[48;2;120;101;104m \033[48;2;160;140;145m \033[48;2;164;147;153m \033[48;2;156;138;147m \033[48;2;175;158;169m \033[48;2;185;164;172m \033[48;2;192;172;181m \033[48;2;173;151;162m \033[48;2;168;147;162m \033[48;2;158;137;152m \033[48;2;143;121;138m \033[48;2;148;128;141m \033[48;2;152;133;152m \033[48;2;152;137;161m \033[48;2;150;138;159m \033[48;2;153;141;163m \033[48;2;157;145;167m \033[48;2;159;146;172m \033[48;2;159;146;172m \033[48;2;156;143;169m \033[48;2;153;137;164m \033[48;2;97;80;102m \033[48;2;69;49;65m \033[48;2;64;47;48m \033[48;2;62;52;48m \033[48;2;58;55;45m \033[48;2;57;53;44m \033[48;2;57;53;44m \033[48;2;57;53;44m \033[48;2;58;50;41m \033[48;2;58;52;40m \033[48;2;56;50;34m \033[48;2;55;52;35m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;52;49;30m \033[48;2;52;49;30m \033[48;2;51;48;29m \033[48;2;51;48;29m \033[48;2;51;48;29m \033[48;2;52;49;30m \033[48;2;52;49;32m \033[48;2;52;49;32m \033[48;2;55;52;35m \033[48;2;57;54;37m \033[48;2;53;50;33m \033[48;2;48;45;28m \033[48;2;51;45;29m \033[48;2;51;48;33m \033[48;2;52;53;39m \033[48;2;54;55;48m \033[48;2;58;57;52m \033[48;2;58;57;52m \033[48;2;60;58;61m \033[48;2;61;59;62m \033[48;2;54;52;55m \033[48;2;53;54;54m \033[48;2;58;58;59m \033[48;2;61;61;61m \033[48;2;60;61;62m \033[48;2;60;60;63m \033[48;2;60;60;63m \033[48;2;60;60;63m \033[48;2;60;60;63m \033[48;2;61;60;63m \033[48;2;69;66;71m \033[48;2;78;69;80m \033[48;2;138;124;141m \033[48;2;170;153;172m \033[48;2;167;152;173m \033[48;2;166;151;176m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[m");
$display("\033[48;2;168;149;171m \033[48;2;168;149;171m \033[48;2;166;148;170m \033[48;2;171;149;172m \033[48;2;141;117;141m \033[48;2;85;53;66m \033[48;2;75;50;53m \033[48;2;71;54;45m \033[48;2;66;57;40m \033[48;2;65;56;39m \033[48;2;65;56;39m \033[48;2;64;57;39m \033[48;2;65;58;40m \033[48;2;70;63;45m \033[48;2;59;52;34m \033[48;2;63;56;38m \033[48;2;59;52;34m \033[48;2;59;52;34m \033[48;2;58;51;33m \033[48;2;56;49;31m \033[48;2;55;50;31m \033[48;2;55;50;31m \033[48;2;55;50;31m \033[48;2;57;52;33m \033[48;2;57;52;30m \033[48;2;57;53;28m \033[48;2;58;53;33m \033[48;2;58;53;33m \033[48;2;59;54;34m \033[48;2;63;54;37m \033[48;2;85;72;57m \033[48;2;107;89;76m \033[48;2;91;74;59m \033[48;2;74;58;42m \033[48;2;73;57;42m \033[48;2;79;61;49m \033[48;2;90;72;65m \033[48;2;93;74;71m \033[48;2;94;75;71m \033[48;2;106;84;83m \033[48;2;119;92;97m \033[48;2;105;77;76m \033[48;2;91;61;62m \033[48;2;89;61;60m \033[48;2;95;76;72m \033[48;2;103;85;80m \033[48;2;114;95;91m \033[48;2;116;98;93m \033[48;2;109;91;89m \033[48;2;101;82;83m \033[48;2;121;105;108m \033[48;2;148;131;137m \033[48;2;166;149;160m \033[48;2;157;141;160m \033[48;2;159;145;167m \033[48;2;143;129;145m \033[48;2;130;112;123m \033[48;2;128;112;122m \033[48;2;116;99;106m \033[48;2;63;54;49m \033[48;2;60;53;47m \033[48;2;55;52;45m \033[48;2;56;52;40m \033[48;2;56;52;40m \033[48;2;55;51;39m \033[48;2;53;52;36m \033[48;2;52;53;35m \033[48;2;50;51;33m \033[48;2;53;50;31m \033[48;2;53;50;31m \033[48;2;52;49;30m \033[48;2;52;50;29m \033[48;2;52;50;29m \033[48;2;52;50;29m \033[48;2;52;49;30m \033[48;2;52;49;30m \033[48;2;54;51;32m \033[48;2;53;50;33m \033[48;2;53;50;33m \033[48;2;53;50;33m \033[48;2;51;50;32m \033[48;2;49;48;30m \033[48;2;47;46;28m \033[48;2;50;47;33m \033[48;2;50;51;37m \033[48;2;49;52;41m \033[48;2;51;56;51m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;179;23;24m \033[48;2;56;57;52m \033[48;2;56;57;52m \033[48;2;56;57;52m \033[48;2;56;57;52m \033[48;2;53;55;47m \033[48;2;54;55;47m \033[48;2;53;54;47m \033[48;2;53;52;48m \033[48;2;57;55;57m \033[48;2;64;62;66m \033[48;2;73;65;74m \033[48;2;98;86;100m \033[48;2;168;154;170m \033[48;2;169;154;175m \033[48;2;167;152;177m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;165;149;175m \033[m");
$display("\033[48;2;169;150;172m \033[48;2;166;147;169m \033[48;2;166;148;170m \033[48;2;173;150;174m \033[48;2;127;104;127m \033[48;2;86;54;68m \033[48;2;72;48;51m \033[48;2;68;52;43m \033[48;2;62;53;36m \033[48;2;61;52;35m \033[48;2;61;52;35m \033[48;2;61;54;37m \033[48;2;66;59;41m \033[48;2;65;58;40m \033[48;2;59;52;34m \033[48;2;58;51;33m \033[48;2;58;51;33m \033[48;2;58;52;33m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;59;53;35m \033[48;2;59;54;35m \033[48;2;60;55;36m \033[48;2;79;74;55m \033[48;2;106;95;84m \033[48;2;112;99;90m \033[48;2;148;134;129m \033[48;2;157;138;133m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;138;119;116m \033[48;2;139;120;116m \033[48;2;140;121;121m \033[48;2;136;118;114m \033[48;2;138;121;112m \033[48;2;140;124;117m \033[48;2;137;122;117m \033[48;2;123;121;121m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;50;50;32m \033[48;2;51;48;29m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;56;47;26m \033[48;2;51;48;29m \033[48;2;51;48;29m \033[48;2;51;48;29m \033[48;2;57;47;31m \033[48;2;57;45;32m \033[48;2;62;51;37m \033[48;2;59;49;35m \033[48;2;49;41;25m \033[48;2;55;46;31m \033[48;2;53;46;33m \033[48;2;54;49;37m \033[48;2;54;51;42m \033[48;2;57;57;52m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;105;44;39m \033[48;2;53;54;49m \033[48;2;50;51;46m \033[48;2;52;53;48m \033[48;2;52;53;47m \033[48;2;52;53;46m \033[48;2;55;56;48m \033[48;2;55;56;49m \033[48;2;57;56;52m \033[48;2;59;56;58m \033[48;2;62;58;62m \033[48;2;69;62;70m \033[48;2;96;85;99m \033[48;2;172;156;174m \033[48;2;170;155;176m \033[48;2;167;152;176m \033[48;2;167;151;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[m");
$display("\033[48;2;167;148;170m \033[48;2;167;148;170m \033[48;2;166;149;167m \033[48;2;174;148;165m \033[48;2;109;81;95m \033[48;2;82;54;61m \033[48;2;67;48;42m \033[48;2;63;51;34m \033[48;2;60;54;31m \033[48;2;60;54;31m \033[48;2;60;54;31m \033[48;2;60;56;30m \033[48;2;66;61;41m \033[48;2;63;58;39m \033[48;2;58;53;34m \033[48;2;57;52;33m \033[48;2;57;52;33m \033[48;2;55;53;32m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;57;53;34m \033[48;2;58;52;38m \033[48;2;58;52;38m \033[48;2;66;60;47m \033[48;2;92;84;71m \033[48;2;91;81;70m \033[48;2;111;96;91m \033[48;2;253;18;19m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;65;52;44m \033[48;2;61;47;37m \033[48;2;62;47;40m \033[48;2;63;49;41m \033[48;2;66;52;44m \033[48;2;66;53;43m \033[48;2;62;59;49m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;52;49;30m \033[48;2;51;48;29m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;56;46;27m \033[48;2;47;48;28m \033[48;2;49;48;28m \033[48;2;49;47;23m \033[48;2;63;51;30m \033[48;2;103;71;56m \033[48;2;143;92;83m \033[48;2;169;107;97m \033[48;2;163;94;92m \033[48;2;159;95;100m \033[48;2;84;43;45m \033[48;2;75;46;49m \033[48;2;68;56;55m \033[48;2;63;59;59m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;31;51;36m \033[48;2;47;47;35m \033[48;2;52;52;42m \033[48;2;55;54;49m \033[48;2;54;53;49m \033[48;2;54;53;49m \033[48;2;51;49;50m \033[48;2;60;55;54m \033[48;2;61;55;55m \033[48;2;61;55;59m \033[48;2;61;54;63m \033[48;2;70;60;71m \033[48;2;123;110;126m \033[48;2;172;157;177m \033[48;2;171;156;177m \033[48;2;170;155;176m \033[48;2;170;155;177m \033[48;2;166;150;176m \033[48;2;166;150;176m \033[m");
$display("\033[48;2;169;151;167m \033[48;2;169;151;167m \033[48;2;165;152;164m \033[48;2;163;142;154m \033[48;2;87;61;74m \033[48;2;75;50;47m \033[48;2;64;51;35m \033[48;2;60;55;27m \033[48;2;59;55;26m \033[48;2;59;55;26m \033[48;2;59;55;26m \033[48;2;59;55;28m \033[48;2;64;59;36m \033[48;2;62;57;37m \033[48;2;58;53;33m \033[48;2;57;52;32m \033[48;2;57;52;32m \033[48;2;55;52;33m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;79;47;30m \033[48;2;55;52;33m \033[48;2;55;52;33m \033[48;2;55;52;33m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;57;54;37m \033[48;2;57;54;37m \033[48;2;68;65;48m \033[48;2;80;74;63m \033[48;2;91;82;75m \033[48;2;114;103;99m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;142;128;126m \033[48;2;154;138;139m \033[48;2;161;145;145m \033[48;2;148;132;133m \033[48;2;144;128;129m \033[48;2;142;126;126m \033[48;2;134;119;119m \033[48;2;137;117;118m \033[48;2;127;109;109m \033[48;2;115;97;96m \033[48;2;102;86;85m \033[48;2;158;43;42m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;55;51;39m \033[48;2;52;49;34m \033[48;2;51;48;29m \033[48;2;50;47;28m \033[48;2;50;47;28m \033[48;2;51;48;29m \033[48;2;51;49;28m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;56;45;26m \033[48;2;44;47;26m \033[48;2;50;48;28m \033[48;2;55;49;27m \033[48;2;61;50;30m \033[48;2;103;75;62m \033[48;2;143;90;84m \033[48;2;142;73;75m \033[48;2;152;74;85m \033[48;2;157;87;97m \033[48;2;140;84;98m \033[48;2;86;44;55m \033[48;2;75;54;55m \033[48;2;60;50;48m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;51;58;50m \033[48;2;55;54;51m \033[48;2;54;53;52m \033[48;2;51;50;47m \033[48;2;54;53;49m \033[48;2;57;56;52m \033[48;2;59;58;54m \033[48;2;57;54;51m \033[48;2;57;51;51m \033[48;2;59;53;57m \033[48;2;65;54;63m \033[48;2;102;90;102m \033[48;2;170;153;173m \033[48;2;175;156;178m \033[48;2;174;155;177m \033[48;2;174;155;177m \033[48;2;174;155;177m \033[48;2;170;155;176m \033[48;2;166;150;176m \033[m");
$display("\033[48;2;167;151;168m \033[48;2;168;151;168m \033[48;2;165;152;166m \033[48;2;156;135;148m \033[48;2;80;54;68m \033[48;2;76;53;47m \033[48;2;67;55;36m \033[48;2;63;58;30m \033[48;2;60;56;28m \033[48;2;59;55;27m \033[48;2;59;55;27m \033[48;2;59;55;29m \033[48;2;62;58;34m \033[48;2;60;56;33m \033[48;2;58;53;33m \033[48;2;57;52;32m \033[48;2;57;52;32m \033[48;2;54;52;32m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;81;49;31m \033[48;2;56;53;34m \033[48;2;55;52;32m \033[48;2;55;53;33m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;55;52;35m \033[48;2;57;54;37m \033[48;2;66;63;46m \033[48;2;94;88;78m \033[48;2;108;98;92m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;162;139;156m \033[48;2;160;123;136m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;64;50;43m \033[48;2;59;47;39m \033[48;2;56;42;34m \033[48;2;53;39;27m \033[48;2;55;41;30m \033[48;2;58;44;33m \033[48;2;59;44;29m \033[48;2;62;47;32m \033[48;2;72;57;43m \033[48;2;72;57;52m \033[48;2;150;35;31m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;54;50;38m \033[48;2;50;46;32m \033[48;2;50;47;29m \033[48;2;49;46;27m \033[48;2;49;47;27m \033[48;2;50;48;26m \033[48;2;51;49;27m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;55;47;27m \033[48;2;44;50;28m \033[48;2;46;51;29m \033[48;2;54;52;29m \033[48;2;63;50;32m \033[48;2;101;74;59m \033[48;2;144;90;83m \033[48;2;135;67;67m \033[48;2;145;69;77m \033[48;2;150;83;92m \033[48;2;154;93;103m \033[48;2;103;53;60m \033[48;2;66;40;38m \033[48;2;50;39;28m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;54;51;42m \033[48;2;57;53;49m \033[48;2;55;51;46m \033[48;2;55;48;44m \033[48;2;54;51;44m \033[48;2;48;47;39m \033[48;2;52;52;47m \033[48;2;56;52;48m \033[48;2;65;58;58m \033[48;2;75;70;74m \033[48;2;112;101;113m \033[48;2;165;153;168m \033[48;2;171;154;173m \033[48;2;173;154;177m \033[48;2;174;155;177m \033[48;2;175;156;178m \033[48;2;175;156;178m \033[48;2;173;155;178m \033[48;2;169;151;177m \033[m");
$display("\033[48;2;165;151;168m \033[48;2;165;151;168m \033[48;2;165;151;168m \033[48;2;162;140;158m \033[48;2;83;57;74m \033[48;2;77;53;50m \033[48;2;68;55;38m \033[48;2;64;57;38m \033[48;2;61;56;34m \033[48;2;58;53;31m \033[48;2;58;53;31m \033[48;2;58;53;34m \033[48;2;61;56;37m \033[48;2;59;54;35m \033[48;2;58;53;33m \033[48;2;57;52;32m \033[48;2;57;52;32m \033[48;2;53;51;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;81;50;29m \033[48;2;57;55;34m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;58;53;34m \033[48;2;55;52;35m \033[48;2;55;52;35m \033[48;2;62;59;42m \033[48;2;68;60;51m \033[48;2;77;65;60m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;154;136;150m \033[48;2;148;131;143m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;190;65;63m \033[48;2;131;120;115m \033[48;2;132;122;119m \033[48;2;135;120;113m \033[48;2;137;122;115m \033[48;2;142;127;120m \033[48;2;140;124;125m \033[48;2;138;121;122m \033[48;2;131;115;115m \033[48;2;124;109;104m \033[48;2;173;62;58m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;53;49;38m \033[48;2;51;47;35m \033[48;2;48;45;28m \033[48;2;48;45;26m \033[48;2;48;46;25m \033[48;2;48;46;22m \033[48;2;50;48;25m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;53;48;27m \033[48;2;45;51;28m \033[48;2;48;53;31m \033[48;2;56;53;30m \033[48;2;60;53;33m \033[48;2;71;52;36m \033[48;2;118;81;70m \033[48;2;130;64;63m \033[48;2;131;59;65m \033[48;2;138;72;80m \033[48;2;141;80;89m \033[48;2;114;62;67m \033[48;2;71;32;33m \033[48;2;57;34;26m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;130;106;99m \033[48;2;154;121;114m \033[48;2;151;114;108m \033[48;2;140;98;95m \033[48;2;86;45;44m \033[48;2;76;45;43m \033[48;2;73;54;53m \033[48;2;71;61;62m \033[48;2;70;63;70m \033[48;2;95;88;102m \033[48;2;165;153;170m \033[48;2;166;153;171m \033[48;2;171;153;175m \033[48;2;172;153;176m \033[48;2;172;153;175m \033[48;2;173;154;176m \033[48;2;173;154;176m \033[48;2;173;153;178m \033[48;2;174;154;179m \033[m");
$display("\033[48;2;166;152;167m \033[48;2;166;152;167m \033[48;2;166;152;169m \033[48;2;166;145;163m \033[48;2;104;76;98m \033[48;2;78;53;56m \033[48;2;68;54;45m \033[48;2;64;58;37m \033[48;2;59;56;37m \033[48;2;56;53;34m \033[48;2;56;53;34m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;32m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;55;52;33m \033[48;2;55;52;33m \033[48;2;56;53;34m \033[48;2;62;59;40m \033[48;2;91;86;73m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;152;139;156m \033[48;2;146;133;147m \033[48;2;140;126;139m \033[48;2;116;107;117m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;70;59;58m \033[48;2;65;52;51m \033[48;2;66;51;42m \033[48;2;62;47;39m \033[48;2;57;42;34m \033[48;2;58;44;30m \033[48;2;53;39;26m \033[48;2;56;42;29m \033[48;2;59;45;32m \033[48;2;140;25;17m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;51;47;36m \033[48;2;48;44;32m \033[48;2;48;45;28m \033[48;2;47;44;25m \033[48;2;47;45;24m \033[48;2;48;46;25m \033[48;2;47;47;23m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;54;48;26m \033[48;2;45;49;26m \033[48;2;48;52;29m \033[48;2;52;51;30m \033[48;2;53;53;28m \033[48;2;53;47;26m \033[48;2;85;57;42m \033[48;2;133;85;81m \033[48;2;131;72;72m \033[48;2;142;76;83m \033[48;2;148;85;94m \033[48;2;143;86;93m \033[48;2;82;37;40m \033[48;2;74;39;37m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;158;116;111m \033[48;2;165;116;110m \033[48;2;170;122;115m \033[48;2;173;124;117m \033[48;2;170;120;115m \033[48;2;128;88;87m \033[48;2;81;55;58m \033[48;2;69;54;59m \033[48;2;66;55;65m \033[48;2;73;61;73m \033[48;2;144;130;145m \033[48;2;173;156;171m \033[48;2;172;153;173m \033[48;2;173;153;176m \033[48;2;173;154;176m \033[48;2;174;155;177m \033[48;2;173;155;177m \033[48;2;170;155;176m \033[48;2;172;157;178m \033[m");
$display("\033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;171;153;174m \033[48;2;129;106;130m \033[48;2;79;52;64m \033[48;2;71;52;48m \033[48;2;64;53;36m \033[48;2;61;55;32m \033[48;2;55;53;31m \033[48;2;54;53;31m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;32m \033[48;2;54;55;28m \033[48;2;51;56;26m \033[48;2;55;53;32m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;52;54;33m \033[48;2;53;53;33m \033[48;2;53;54;33m \033[48;2;55;56;35m \033[48;2;203;23;17m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;240;50;54m \033[48;2;162;144;161m \033[48;2;160;143;157m \033[48;2;136;119;129m \033[48;2;94;80;78m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;125;117;109m \033[48;2;128;117;112m \033[48;2;135;124;119m \033[48;2;135;122;117m \033[48;2;137;121;123m \033[48;2;137;121;120m \033[48;2;136;120;121m \033[48;2;134;119;117m \033[48;2;175;65;63m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;47;43;31m \033[48;2;47;44;29m \033[48;2;48;45;26m \033[48;2;47;45;24m \033[48;2;47;45;24m \033[48;2;47;45;24m \033[48;2;45;46;18m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;54;43;24m \033[48;2;47;45;24m \033[48;2;49;47;26m \033[48;2;52;50;29m \033[48;2;50;50;29m \033[48;2;56;53;33m \033[48;2;75;54;41m \033[48;2;136;94;93m \033[48;2;127;69;72m \033[48;2;138;71;80m \033[48;2;159;96;103m \033[48;2;157;100;106m \033[48;2;140;90;94m \033[48;2;108;65;63m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;169;120;109m \033[48;2;161;105;91m \033[48;2;145;89;74m \033[48;2;128;75;62m \033[48;2;117;71;63m \033[48;2;102;65;57m \033[48;2;79;56;51m \033[48;2;61;49;47m \033[48;2;62;52;53m \033[48;2;75;64;70m \033[48;2;134;120;129m \033[48;2;172;154;168m \033[48;2;172;153;172m \033[48;2;172;153;174m \033[48;2;172;153;175m \033[48;2;173;154;176m \033[48;2;172;154;176m \033[48;2;170;155;176m \033[48;2;171;156;177m \033[m");
$display("\033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;170;152;171m \033[48;2;150;128;151m \033[48;2;85;56;74m \033[48;2;70;50;51m \033[48;2;63;51;40m \033[48;2;60;54;32m \033[48;2;56;53;30m \033[48;2;54;54;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;55;53;32m \033[48;2;52;55;28m \033[48;2;51;56;26m \033[48;2;55;53;32m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;77;49;27m \033[48;2;52;54;30m \033[48;2;52;54;30m \033[48;2;52;54;30m \033[48;2;52;54;30m \033[48;2;52;54;30m \033[48;2;52;54;30m \033[48;2;52;55;28m \033[48;2;52;54;30m \033[48;2;50;52;31m \033[48;2;52;54;33m \033[48;2;52;54;33m \033[48;2;56;58;37m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;114;83;74m \033[48;2;158;123;112m \033[48;2;144;112;102m \033[48;2;129;94;96m \033[48;2;125;91;95m \033[48;2;127;94;92m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;77;69;62m \033[48;2;72;62;53m \033[48;2;69;59;50m \033[48;2;63;53;43m \033[48;2;62;49;38m \033[48;2;60;45;35m \033[48;2;54;40;28m \033[48;2;51;37;26m \033[48;2;134;18;10m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;47;43;31m \033[48;2;47;44;29m \033[48;2;47;44;25m \033[48;2;47;45;24m \033[48;2;47;45;24m \033[48;2;47;45;24m \033[48;2;44;46;18m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;54;43;24m \033[48;2;47;45;24m \033[48;2;49;47;26m \033[48;2;51;49;28m \033[48;2;50;49;29m \033[48;2;50;45;26m \033[48;2;70;50;36m \033[48;2;128;92;89m \033[48;2;122;71;75m \033[48;2;132;71;78m \033[48;2;133;70;79m \033[48;2;140;83;89m \033[48;2;136;83;88m \033[48;2;139;91;92m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;136;81;76m \033[48;2;130;74;71m \033[48;2;115;64;59m \033[48;2;112;64;60m \033[48;2;94;55;54m \033[48;2;78;52;52m \033[48;2;68;54;58m \033[48;2;75;64;69m \033[48;2;75;64;72m \033[48;2;132;120;132m \033[48;2;178;162;173m \033[48;2;173;155;168m \033[48;2;172;153;172m \033[48;2;172;153;174m \033[48;2;172;153;175m \033[48;2;171;152;174m \033[48;2;173;155;177m \033[48;2;171;156;177m \033[48;2;171;156;177m \033[m");
$display("\033[48;2;166;152;167m \033[48;2;166;152;167m \033[48;2;167;153;169m \033[48;2;169;151;168m \033[48;2;163;142;159m \033[48;2;92;65;82m \033[48;2;73;47;55m \033[48;2;65;50;39m \033[48;2;59;52;33m \033[48;2;56;54;29m \033[48;2;55;55;27m \033[48;2;58;53;31m \033[48;2;58;53;31m \033[48;2;57;52;30m \033[48;2;53;51;30m \033[48;2;50;52;30m \033[48;2;49;53;30m \033[48;2;53;51;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;79;47;30m \033[48;2;53;50;31m \033[48;2;55;52;33m \033[48;2;55;52;33m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;53;50;31m \033[48;2;52;49;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;122;108;99m \033[48;2;122;108;98m \033[48;2;127;113;105m \033[48;2;127;113;104m \033[48;2;133;118;108m \033[48;2;131;117;107m \033[48;2;129;118;109m \033[48;2;175;68;61m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;46;43;28m \033[48;2;49;46;26m \033[48;2;47;45;24m \033[48;2;47;45;22m \033[48;2;47;45;22m \033[48;2;46;44;21m \033[48;2;46;44;21m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;53;43;20m \033[48;2;49;44;24m \033[48;2;47;45;24m \033[48;2;49;48;27m \033[48;2;44;47;22m \033[48;2;56;51;29m \033[48;2;72;58;39m \033[48;2;121;90;81m \033[48;2;127;77;78m \033[48;2;131;72;78m \033[48;2;130;77;81m \033[48;2;129;77;81m \033[48;2;136;84;88m \033[48;2;134;82;81m \033[48;2;136;85;82m \033[48;2;139;88;85m \033[48;2;167;116;113m \033[48;2;173;122;119m \033[48;2;159;107;113m \033[48;2;151;100;111m \033[48;2;132;84;100m \033[48;2;87;44;65m \033[48;2;81;51;65m \033[48;2;72;54;63m \033[48;2;66;61;61m \033[48;2;66;61;62m \033[48;2;91;85;92m \033[48;2;166;151;163m \033[48;2;172;154;170m \033[48;2;174;156;172m \033[48;2;174;156;172m \033[48;2;173;154;173m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;172;153;175m \033[48;2;170;155;176m \033[48;2;171;156;177m \033[m");
$display("\033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;167;153;166m \033[48;2;171;153;167m \033[48;2;161;140;155m \033[48;2;90;67;78m \033[48;2;75;53;51m \033[48;2;62;51;33m \033[48;2;60;53;34m \033[48;2;57;54;33m \033[48;2;55;54;33m \033[48;2;58;53;31m \033[48;2;58;53;31m \033[48;2;57;52;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;77;49;30m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;53;51;30m \033[48;2;50;52;30m \033[48;2;43;54;31m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;135;125;119m \033[48;2;98;84;82m \033[48;2;125;107;109m \033[48;2;121;107;105m \033[48;2;126;112;107m \033[48;2;129;115;108m \033[48;2;124;109;105m \033[48;2;121;107;103m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;152;55;48m \033[48;2;85;71;61m \033[48;2;74;58;50m \033[48;2;72;57;53m \033[48;2;65;50;46m \033[48;2;60;44;39m \033[48;2;56;41;33m \033[48;2;138;22;17m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;42;43;27m \033[48;2;42;44;23m \033[48;2;42;44;22m \033[48;2;43;45;21m \033[48;2;43;45;21m \033[48;2;43;45;21m \033[48;2;43;45;23m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;53;42;18m \033[48;2;42;42;13m \033[48;2;45;43;18m \033[48;2;48;46;24m \033[48;2;49;49;29m \033[48;2;52;50;31m \033[48;2;71;53;39m \033[48;2;124;88;81m \033[48;2;122;79;73m \033[48;2;127;74;71m \033[48;2;151;97;95m \033[48;2;142;91;88m \033[48;2;139;88;86m \033[48;2;139;82;81m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;145;104;105m \033[48;2;152;103;108m \033[48;2;149;104;114m \033[48;2;120;79;100m \033[48;2;78;48;65m \033[48;2;70;53;60m \033[48;2;63;55;55m \033[48;2;59;58;53m \033[48;2;64;61;56m \033[48;2;71;69;63m \033[48;2;124;112;113m \033[48;2;170;152;162m \033[48;2;175;157;175m \033[48;2;174;156;175m \033[48;2;171;156;175m \033[48;2;170;155;176m \033[48;2;170;155;176m \033[48;2;170;156;173m \033[48;2;171;157;174m \033[m");
$display("\033[48;2;167;153;168m \033[48;2;167;153;168m \033[48;2;167;153;166m \033[48;2;170;152;166m \033[48;2;157;136;151m \033[48;2;84;61;72m \033[48;2;70;50;48m \033[48;2;62;50;34m \033[48;2;60;53;34m \033[48;2;57;54;33m \033[48;2;55;54;33m \033[48;2;58;53;31m \033[48;2;58;53;31m \033[48;2;57;52;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;77;49;30m \033[48;2;55;53;32m \033[48;2;54;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;51;52;30m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;57;50;32m \033[48;2;112;101;95m \033[48;2;97;82;79m \033[48;2;121;102;104m \033[48;2;68;52;51m \033[48;2;62;47;42m \033[48;2;66;51;44m \033[48;2;73;59;48m \033[48;2;73;59;50m \033[48;2;242;6;5m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;115;102;87m \033[48;2;113;114;97m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;42;44;20m \033[48;2;43;45;23m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;124;71;69m \033[48;2;145;95;92m \033[48;2;155;104;102m \033[48;2;210;40;41m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;135;85;95m \033[48;2;134;88;98m \033[48;2;118;82;86m \033[48;2;83;56;56m \033[48;2;75;60;56m \033[48;2;68;59;57m \033[48;2;61;60;60m \033[48;2;66;62;63m \033[48;2;59;53;55m \033[48;2;58;48;47m \033[48;2;78;67;68m \033[48;2;134;123;132m \033[48;2;168;154;170m \033[48;2;167;153;171m \033[48;2;170;155;176m \033[48;2;170;155;178m \033[48;2;168;153;177m \033[48;2;169;154;177m \033[m");
$display("\033[48;2;168;154;169m \033[48;2;168;154;169m \033[48;2;170;153;169m \033[48;2;176;154;172m \033[48;2;152;129;147m \033[48;2;83;52;63m \033[48;2;68;44;44m \033[48;2;61;49;37m \033[48;2;60;53;34m \033[48;2;60;53;34m \033[48;2;60;53;34m \033[48;2;58;53;33m \033[48;2;56;51;31m \033[48;2;56;51;31m \033[48;2;54;52;31m \033[48;2;54;52;31m \033[48;2;54;52;31m \033[48;2;51;53;29m \033[48;2;49;52;28m \033[48;2;50;53;28m \033[48;2;51;54;29m \033[48;2;51;54;29m \033[48;2;51;53;29m \033[48;2;51;53;29m \033[48;2;49;51;27m \033[48;2;49;51;27m \033[48;2;52;50;29m \033[48;2;52;50;29m \033[48;2;52;50;29m \033[48;2;53;51;28m \033[48;2;54;52;29m \033[48;2;52;50;27m \033[48;2;52;51;23m \033[48;2;53;52;27m \033[48;2;54;53;31m \033[48;2;56;52;33m \033[48;2;77;72;57m \033[48;2;125;119;107m \033[48;2;131;120;114m \033[48;2;110;96;94m \033[48;2;123;102;104m \033[48;2;132;114;110m \033[48;2;133;115;111m \033[48;2;135;117;113m \033[48;2;131;116;111m \033[48;2;129;114;112m \033[48;2;125;109;110m \033[48;2;121;107;109m \033[48;2;117;103;103m \033[48;2;111;97;98m \033[48;2;104;92;84m \033[48;2;97;83;77m \033[48;2;88;73;69m \033[48;2;77;64;55m \033[48;2;77;64;54m \033[48;2;69;57;47m \033[48;2;64;51;41m \033[48;2;54;41;31m \033[48;2;54;40;30m \033[48;2;52;40;30m \033[48;2;56;50;39m \033[48;2;58;52;40m \033[48;2;46;46;31m \033[48;2;40;42;21m \033[48;2;39;41;19m \033[48;2;40;43;18m \033[48;2;40;43;18m \033[48;2;40;42;18m \033[48;2;40;43;17m \033[48;2;40;44;17m \033[48;2;40;44;17m \033[48;2;40;44;17m \033[48;2;40;44;17m \033[48;2;40;42;16m \033[48;2;43;43;14m \033[48;2;43;43;14m \033[48;2;42;41;13m \033[48;2;44;44;15m \033[48;2;55;54;29m \033[48;2;63;48;30m \033[48;2;96;61;53m \033[48;2;122;79;75m \033[48;2;121;69;67m \033[48;2;131;71;70m \033[48;2;140;80;78m \033[48;2;149;90;92m \033[48;2;153;93;100m \033[48;2;155;99;106m \033[48;2;255;0;0m \033[48;2;255;0;0m \033[48;2;160;113;119m \033[48;2;154;107;113m \033[48;2;155;110;117m \033[48;2;129;88;93m \033[48;2;80;47;52m \033[48;2;71;49;49m \033[48;2;64;51;50m \033[48;2;62;58;55m \033[48;2;60;60;62m \033[48;2;60;60;62m \033[48;2;61;61;63m \033[48;2;61;62;64m \033[48;2;62;61;63m \033[48;2;69;63;67m \033[48;2;104;96;101m \033[48;2;160;147;158m \033[48;2;171;158;175m \033[48;2;171;157;181m \033[48;2;171;155;179m \033[48;2;171;156;177m \033[m");
$display("\033[48;2;170;152;168m \033[48;2;170;152;168m \033[48;2;169;153;166m \033[48;2;175;153;168m \033[48;2;151;128;144m \033[48;2;83;53;65m \033[48;2;75;50;52m \033[48;2;65;53;43m \033[48;2;60;53;35m \033[48;2;60;53;35m \033[48;2;60;53;35m \033[48;2;57;52;32m \033[48;2;55;50;30m \033[48;2;55;50;30m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;53;51;28m \033[48;2;50;52;28m \033[48;2;52;54;30m \033[48;2;49;51;27m \033[48;2;54;52;31m \033[48;2;52;50;29m \033[48;2;51;49;28m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;47;49;27m \033[48;2;49;47;28m \033[48;2;56;50;34m \033[48;2;112;102;95m \033[48;2;108;92;91m \033[48;2;108;87;89m \033[48;2;63;45;38m \033[48;2;61;44;35m \033[48;2;64;48;35m \033[48;2;66;53;36m \033[48;2;71;58;41m \033[48;2;72;59;42m \033[48;2;79;67;51m \033[48;2;84;71;55m \033[48;2;93;81;65m \033[48;2;100;87;71m \033[48;2;102;89;73m \033[48;2;113;100;84m \033[48;2;120;106;93m \033[48;2;123;109;98m \033[48;2;126;112;102m \033[48;2;127;110;101m \033[48;2;120;103;94m \033[48;2;115;98;90m \033[48;2;108;92;79m \033[48;2;89;75;61m \033[48;2;62;50;40m \033[48;2;55;50;37m \033[48;2;45;41;27m \033[48;2;39;41;20m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;38;43;13m \033[48;2;41;41;13m \033[48;2;45;37;11m \033[48;2;63;57;38m \033[48;2;80;64;48m \033[48;2;90;57;48m \033[48;2;96;50;43m \033[48;2;126;76;72m \033[48;2;122;67;67m \033[48;2;127;70;71m \033[48;2;129;72;73m \033[48;2;142;82;86m \033[48;2;172;117;121m \033[48;2;148;96;100m \033[48;2;144;92;96m \033[48;2;152;101;106m \033[48;2;147;101;104m \033[48;2;153;108;111m \033[48;2;147;105;107m \033[48;2;129;87;89m \033[48;2;77;48;49m \033[48;2;62;48;45m \033[48;2;54;49;38m \033[48;2;57;59;47m \033[48;2;58;59;53m \033[48;2;58;59;53m \033[48;2;60;59;60m \033[48;2;61;61;60m \033[48;2;61;61;61m \033[48;2;61;60;65m \033[48;2;64;61;67m \033[48;2;98;92;98m \033[48;2;160;149;158m \033[48;2;168;155;171m \033[48;2;167;154;174m \033[48;2;168;155;175m \033[m");
$display("\033[48;2;172;154;170m \033[48;2;172;154;170m \033[48;2;171;155;168m \033[48;2;173;152;167m \033[48;2;155;132;148m \033[48;2;91;60;73m \033[48;2;76;50;53m \033[48;2;63;51;41m \033[48;2;60;53;35m \033[48;2;60;53;35m \033[48;2;60;53;35m \033[48;2;57;52;32m \033[48;2;56;51;31m \033[48;2;57;52;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;32m \033[48;2;55;53;30m \033[48;2;55;53;30m \033[48;2;53;51;28m \033[48;2;50;52;28m \033[48;2;50;52;28m \033[48;2;50;52;28m \033[48;2;54;52;31m \033[48;2;52;50;29m \033[48;2;51;49;28m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;51;49;26m \033[48;2;48;50;27m \033[48;2;52;50;30m \033[48;2;105;99;83m \033[48;2;125;116;109m \033[48;2;114;99;97m \033[48;2;113;93;96m \033[48;2;130;111;117m \033[48;2;134;115;119m \033[48;2;139;121;120m \033[48;2;137;122;118m \033[48;2;129;114;110m \033[48;2;128;113;109m \033[48;2;123;110;102m \033[48;2;122;106;99m \033[48;2;114;100;95m \033[48;2;113;98;91m \033[48;2;106;91;84m \033[48;2;92;78;72m \033[48;2;86;71;62m \033[48;2;79;65;55m \033[48;2;73;58;48m \033[48;2;70;54;40m \033[48;2;70;54;40m \033[48;2;60;44;29m \033[48;2;61;45;26m \033[48;2;59;46;30m \033[48;2;56;45;30m \033[48;2;54;48;36m \033[48;2;54;50;36m \033[48;2;43;44;23m \033[48;2;38;41;12m \033[48;2;38;41;12m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;38;43;13m \033[48;2;41;41;13m \033[48;2;45;38;13m \033[48;2;83;58;42m \033[48;2;127;92;76m \033[48;2;140;91;81m \033[48;2;143;81;79m \033[48;2;147;86;85m \033[48;2;152;95;97m \033[48;2;146;95;95m \033[48;2;150;99;98m \033[48;2;164;113;112m \033[48;2;178;127;131m \033[48;2;174;122;126m \033[48;2;151;99;103m \033[48;2;141;91;96m \033[48;2;143;97;99m \033[48;2;146;101;104m \033[48;2;135;92;98m \033[48;2;107;64;74m \033[48;2;84;51;59m \033[48;2;72;56;62m \033[48;2;56;50;42m \033[48;2;42;43;28m \033[48;2;40;43;25m \033[48;2;42;46;28m \033[48;2;47;49;37m \033[48;2;56;57;48m \033[48;2;57;58;52m \033[48;2;60;60;58m \033[48;2;63;64;65m \033[48;2;66;65;70m \033[48;2;106;102;108m \033[48;2;163;153;168m \033[48;2;165;152;172m \033[48;2;167;154;174m \033[m");
$display("\033[48;2;170;156;171m \033[48;2;170;156;171m \033[48;2;173;157;170m \033[48;2;173;153;167m \033[48;2;163;140;156m \033[48;2;106;78;93m \033[48;2;76;49;56m \033[48;2;68;51;44m \033[48;2;63;56;38m \033[48;2;63;56;38m \033[48;2;59;52;34m \033[48;2;56;51;31m \033[48;2;54;49;24m \033[48;2;53;49;22m \033[48;2;53;51;30m \033[48;2;52;50;29m \033[48;2;52;50;29m \033[48;2;52;50;25m \033[48;2;52;50;26m \033[48;2;54;52;26m \033[48;2;51;53;29m \033[48;2;49;51;27m \033[48;2;49;51;27m \033[48;2;48;50;26m \033[48;2;48;50;26m \033[48;2;47;49;25m \033[48;2;47;50;21m \033[48;2;47;50;21m \033[48;2;47;50;21m \033[48;2;47;50;21m \033[48;2;47;50;21m \033[48;2;47;50;21m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;50;23m \033[48;2;51;50;27m \033[48;2;58;53;35m \033[48;2;112;102;95m \033[48;2;107;91;95m \033[48;2;93;73;75m \033[48;2;63;46;40m \033[48;2;59;42;32m \033[48;2;59;43;30m \033[48;2;54;41;24m \033[48;2;58;45;28m \033[48;2;59;47;30m \033[48;2;62;48;35m \033[48;2;70;56;43m \033[48;2;74;60;47m \033[48;2;82;68;57m \033[48;2;90;76;64m \033[48;2;95;81;70m \033[48;2;103;89;78m \033[48;2;114;100;87m \033[48;2;119;105;93m \033[48;2;121;107;97m \033[48;2;106;92;81m \033[48;2;101;89;73m \033[48;2;96;85;66m \033[48;2;95;82;64m \033[48;2;89;76;58m \033[48;2;57;53;34m \033[48;2;51;48;29m \033[48;2;46;47;26m \033[48;2;38;40;16m \033[48;2;38;41;14m \033[48;2;38;41;10m \033[48;2;38;41;12m \033[48;2;38;41;12m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;39;42;13m \033[48;2;36;41;11m \033[48;2;43;38;11m \033[48;2;55;41;23m \033[48;2;103;63;56m \033[48;2;138;86;86m \033[48;2;149;84;92m \033[48;2;146;84;94m \033[48;2;158;99;110m \033[48;2;154;99;107m \033[48;2;152;100;104m \033[48;2;164;112;114m \033[48;2;163;114;117m \033[48;2;165;116;119m \033[48;2;154;105;108m \033[48;2;152;105;110m \033[48;2;154;109;114m \033[48;2;150;108;112m \033[48;2;135;96;95m \033[48;2;130;89;91m \033[48;2;80;51;52m \033[48;2;70;56;56m \033[48;2;65;54;52m \033[48;2;62;58;49m \033[48;2;59;59;49m \033[48;2;55;57;49m \033[48;2;54;55;51m \033[48;2;54;56;50m \033[48;2;58;59;54m \033[48;2;61;61;61m \033[48;2;62;62;62m \033[48;2;62;60;66m \033[48;2;68;67;73m \033[48;2;118;112;125m \033[48;2;162;149;169m \033[48;2;164;151;171m \033[m");
$display("\033[48;2;170;156;171m \033[48;2;170;156;171m \033[48;2;167;153;168m \033[48;2;170;152;168m \033[48;2;166;145;162m \033[48;2;130;102;119m \033[48;2;78;51;58m \033[48;2;69;53;49m \033[48;2;64;55;40m \033[48;2;62;55;37m \033[48;2;57;54;32m \033[48;2;54;49;30m \033[48;2;52;47;24m \033[48;2;52;48;21m \033[48;2;52;51;22m \033[48;2;53;51;28m \033[48;2;53;51;30m \033[48;2;53;51;28m \033[48;2;53;51;28m \033[48;2;53;51;28m \033[48;2;50;52;28m \033[48;2;49;51;27m \033[48;2;49;51;27m \033[48;2;48;52;27m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;46;50;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;46;49;19m \033[48;2;51;51;24m \033[48;2;80;75;55m \033[48;2;119;109;98m \033[48;2;111;98;94m \033[48;2;98;80;78m \033[48;2;126;111;108m \033[48;2;129;114;110m \033[48;2;133;119;109m \033[48;2;134;120;111m \033[48;2;132;118;110m \033[48;2;128;114;105m \033[48;2;124;110;103m \033[48;2;123;108;102m \033[48;2;116;102;94m \033[48;2;110;95;88m \033[48;2;108;93;86m \033[48;2;91;77;70m \033[48;2;84;71;61m \033[48;2;76;62;52m \033[48;2;60;47;37m \033[48;2;56;44;23m \033[48;2;52;39;20m \033[48;2;55;44;24m \033[48;2;61;49;29m \033[48;2;61;49;30m \033[48;2;55;43;24m \033[48;2;54;46;26m \033[48;2;51;46;27m \033[48;2;49;46;30m \033[48;2;42;44;22m \033[48;2;33;35;13m \033[48;2;37;40;12m \033[48;2;38;43;11m \033[48;2;38;43;11m \033[48;2;38;43;11m \033[48;2;38;43;11m \033[48;2;38;43;11m \033[48;2;37;42;10m \033[48;2;37;42;12m \033[48;2;37;38;10m \033[48;2;39;37;9m \033[48;2;41;36;3m \033[48;2;52;34;9m \033[48;2;81;38;29m \033[48;2;104;51;48m \033[48;2;115;61;61m \033[48;2;128;72;74m \033[48;2;148;97;96m \033[48;2;147;95;94m \033[48;2;143;92;93m \033[48;2;138;88;87m \033[48;2;144;96;95m \033[48;2;139;94;91m \033[48;2;133;92;93m \033[48;2;136;96;97m \033[48;2;137;97;98m \033[48;2;135;96;96m \033[48;2;120;80;76m \033[48;2;91;62;52m \033[48;2;68;54;41m \033[48;2;63;51;48m \033[48;2;64;55;58m \033[48;2;62;58;55m \033[48;2;60;59;57m \033[48;2;58;59;62m \033[48;2;55;56;59m \033[48;2;53;53;55m \033[48;2;53;53;55m \033[48;2;54;54;58m \033[48;2;56;57;62m \033[48;2;61;62;67m \033[48;2;70;71;77m \033[48;2;125;122;133m \033[48;2;160;151;167m \033[m");
$display("\033[48;2;170;156;171m \033[48;2;170;156;171m \033[48;2;168;154;169m \033[48;2;170;152;168m \033[48;2;168;147;164m \033[48;2;145;119;136m \033[48;2;78;53;63m \033[48;2;74;56;55m \033[48;2;62;53;38m \033[48;2;59;52;34m \033[48;2;56;52;31m \033[48;2;53;49;30m \033[48;2;50;46;21m \033[48;2;49;46;19m \033[48;2;50;49;21m \033[48;2;53;51;28m \033[48;2;53;51;30m \033[48;2;53;51;29m \033[48;2;53;51;29m \033[48;2;53;51;29m \033[48;2;49;51;27m \033[48;2;48;50;26m \033[48;2;49;51;27m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;46;50;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;46;50;21m \033[48;2;48;48;23m \033[48;2;62;57;36m \033[48;2;112;103;93m \033[48;2;105;91;89m \033[48;2;74;57;54m \033[48;2;62;47;40m \033[48;2;56;43;32m \033[48;2;52;39;28m \033[48;2;51;37;26m \033[48;2;55;41;27m \033[48;2;56;42;31m \033[48;2;57;44;27m \033[48;2;59;46;30m \033[48;2;60;47;29m \033[48;2;67;54;37m \033[48;2;69;55;38m \033[48;2;82;69;52m \033[48;2;93;77;64m \033[48;2;104;90;77m \033[48;2;122;107;94m \033[48;2;120;106;94m \033[48;2;130;115;104m \033[48;2;119;105;93m \033[48;2;109;95;79m \033[48;2;95;83;64m \033[48;2;80;65;49m \033[48;2;72;58;42m \033[48;2;61;48;34m \033[48;2;53;43;29m \033[48;2;51;48;34m \033[48;2;39;39;21m \033[48;2;38;40;18m \033[48;2;37;42;12m \033[48;2;37;42;13m \033[48;2;37;42;10m \033[48;2;37;42;10m \033[48;2;37;42;10m \033[48;2;37;42;12m \033[48;2;34;43;13m \033[48;2;36;42;13m \033[48;2;36;39;11m \033[48;2;33;40;9m \033[48;2;35;40;8m \033[48;2;37;42;9m \033[48;2;44;40;9m \033[48;2;47;35;9m \033[48;2;71;43;24m \033[48;2;86;44;32m \033[48;2;119;74;62m \033[48;2;121;73;63m \033[48;2;119;69;66m \033[48;2;120;71;69m \033[48;2;126;82;78m \033[48;2;130;88;90m \033[48;2;132;92;93m \033[48;2;130;90;91m \033[48;2;121;80;78m \033[48;2;101;63;55m \033[48;2;94;64;48m \033[48;2;64;49;37m \033[48;2;64;54;49m \033[48;2;64;55;56m \033[48;2;61;58;55m \033[48;2;57;57;55m \033[48;2;57;58;60m \033[48;2;57;59;62m \033[48;2;56;58;59m \033[48;2;52;52;55m \033[48;2;50;52;56m \033[48;2;55;57;62m \033[48;2;61;63;68m \033[48;2;62;64;69m \033[48;2;67;66;76m \033[48;2;132;122;136m \033[m");
$display("\033[48;2;171;159;173m \033[48;2;169;157;171m \033[48;2;169;155;170m \033[48;2;171;153;169m \033[48;2;167;146;163m \033[48;2;158;133;148m \033[48;2;86;63;72m \033[48;2;74;52;56m \033[48;2;60;51;36m \033[48;2;58;51;33m \033[48;2;53;50;28m \033[48;2;50;48;27m \033[48;2;48;46;22m \033[48;2;48;47;19m \033[48;2;49;48;20m \033[48;2;52;50;26m \033[48;2;52;50;29m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;53;51;30m \033[48;2;49;51;27m \033[48;2;49;51;27m \033[48;2;49;51;27m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;47;51;26m \033[48;2;46;50;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;47;49;25m \033[48;2;50;50;25m \033[48;2;69;63;42m \033[48;2;117;109;98m \033[48;2;108;97;92m \033[48;2;97;82;79m \033[48;2;120;105;98m \033[48;2;121;106;99m \033[48;2;123;109;101m \033[48;2;130;115;108m \033[48;2;133;118;111m \033[48;2;137;122;115m \033[48;2;136;121;117m \033[48;2;131;116;111m \033[48;2;131;116;111m \033[48;2;127;110;104m \033[48;2;122;105;98m \033[48;2;116;99;92m \033[48;2;109;92;84m \033[48;2;99;82;74m \033[48;2;82;65;57m \033[48;2;77;60;50m \033[48;2;63;46;36m \033[48;2;63;45;36m \033[48;2;53;37;22m \033[48;2;56;40;25m \033[48;2;64;48;33m \033[48;2;71;57;44m \033[48;2;89;75;62m \033[48;2;94;80;67m \033[48;2;69;58;45m \033[48;2;53;45;28m \033[48;2;51;48;28m \033[48;2;41;44;20m \033[48;2;38;42;15m \033[48;2;37;42;10m \033[48;2;36;43;10m \033[48;2;36;43;11m \033[48;2;36;42;15m \033[48;2;37;41;16m \033[48;2;35;39;14m \033[48;2;34;38;13m \033[48;2;36;41;10m \033[48;2;36;41;9m \033[48;2;36;41;9m \033[48;2;33;43;11m \033[48;2;33;42;11m \033[48;2;39;43;14m \033[48;2;53;50;23m \033[48;2;62;48;25m \033[48;2;70;44;23m \033[48;2;81;58;34m \033[48;2;86;61;37m \033[48;2;89;60;39m \033[48;2;91;65;44m \033[48;2;91;66;44m \033[48;2;81;56;34m \033[48;2;61;40;16m \033[48;2;54;33;4m \033[48;2;48;33;8m \033[48;2;54;49;33m \033[48;2;61;57;45m \033[48;2;58;57;52m \033[48;2;58;59;54m \033[48;2;58;58;56m \033[48;2;58;58;60m \033[48;2;57;58;63m \033[48;2;57;58;63m \033[48;2;58;59;64m \033[48;2;54;57;62m \033[48;2;54;57;62m \033[48;2;57;60;65m \033[48;2;61;64;69m \033[48;2;63;64;69m \033[48;2;73;70;77m \033[m");
$display ("-----------------------------------------------------------------------------------------------------");
$display ("                          Never Gonna Give You Up! Never Gonna Let You Down!                         ");
$display ("-----------------------------------------------------------------------------------------------------");
end endtask

endmodule

